
module Register64bit ( clk, rst, in, out );
  input [63:0] in;
  output [63:0] out;
  input clk, rst;
  wire   n2;

  DFFR_X1 out_reg_32_ ( .D(in[32]), .CK(clk), .RN(n2), .Q(out[32]) );
  DFFR_X1 out_reg_63_ ( .D(in[63]), .CK(clk), .RN(n2), .Q(out[63]) );
  DFFR_X1 out_reg_62_ ( .D(in[62]), .CK(clk), .RN(n2), .Q(out[62]) );
  DFFR_X1 out_reg_61_ ( .D(in[61]), .CK(clk), .RN(n2), .Q(out[61]) );
  DFFR_X1 out_reg_60_ ( .D(in[60]), .CK(clk), .RN(n2), .Q(out[60]) );
  DFFR_X1 out_reg_59_ ( .D(in[59]), .CK(clk), .RN(n2), .Q(out[59]) );
  DFFR_X1 out_reg_58_ ( .D(in[58]), .CK(clk), .RN(n2), .Q(out[58]) );
  DFFR_X1 out_reg_57_ ( .D(in[57]), .CK(clk), .RN(n2), .Q(out[57]) );
  DFFR_X1 out_reg_56_ ( .D(in[56]), .CK(clk), .RN(n2), .Q(out[56]) );
  DFFR_X1 out_reg_55_ ( .D(in[55]), .CK(clk), .RN(n2), .Q(out[55]) );
  DFFR_X1 out_reg_54_ ( .D(in[54]), .CK(clk), .RN(n2), .Q(out[54]) );
  DFFR_X1 out_reg_53_ ( .D(in[53]), .CK(clk), .RN(n2), .Q(out[53]) );
  DFFR_X1 out_reg_52_ ( .D(in[52]), .CK(clk), .RN(n2), .Q(out[52]) );
  DFFR_X1 out_reg_51_ ( .D(in[51]), .CK(clk), .RN(n2), .Q(out[51]) );
  DFFR_X1 out_reg_50_ ( .D(in[50]), .CK(clk), .RN(n2), .Q(out[50]) );
  DFFR_X1 out_reg_49_ ( .D(in[49]), .CK(clk), .RN(n2), .Q(out[49]) );
  DFFR_X1 out_reg_48_ ( .D(in[48]), .CK(clk), .RN(n2), .Q(out[48]) );
  DFFR_X1 out_reg_47_ ( .D(in[47]), .CK(clk), .RN(n2), .Q(out[47]) );
  DFFR_X1 out_reg_46_ ( .D(in[46]), .CK(clk), .RN(n2), .Q(out[46]) );
  DFFR_X1 out_reg_45_ ( .D(in[45]), .CK(clk), .RN(n2), .Q(out[45]) );
  DFFR_X1 out_reg_44_ ( .D(in[44]), .CK(clk), .RN(n2), .Q(out[44]) );
  DFFR_X1 out_reg_43_ ( .D(in[43]), .CK(clk), .RN(n2), .Q(out[43]) );
  DFFR_X1 out_reg_42_ ( .D(in[42]), .CK(clk), .RN(n2), .Q(out[42]) );
  DFFR_X1 out_reg_41_ ( .D(in[41]), .CK(clk), .RN(n2), .Q(out[41]) );
  DFFR_X1 out_reg_40_ ( .D(in[40]), .CK(clk), .RN(n2), .Q(out[40]) );
  DFFR_X1 out_reg_39_ ( .D(in[39]), .CK(clk), .RN(n2), .Q(out[39]) );
  DFFR_X1 out_reg_38_ ( .D(in[38]), .CK(clk), .RN(n2), .Q(out[38]) );
  DFFR_X1 out_reg_37_ ( .D(in[37]), .CK(clk), .RN(n2), .Q(out[37]) );
  DFFR_X1 out_reg_36_ ( .D(in[36]), .CK(clk), .RN(n2), .Q(out[36]) );
  DFFR_X1 out_reg_35_ ( .D(in[35]), .CK(clk), .RN(n2), .Q(out[35]) );
  DFFR_X1 out_reg_34_ ( .D(in[34]), .CK(clk), .RN(n2), .Q(out[34]) );
  DFFR_X1 out_reg_33_ ( .D(in[33]), .CK(clk), .RN(n2), .Q(out[33]) );
  DFFR_X1 out_reg_31_ ( .D(in[31]), .CK(clk), .RN(n2), .Q(out[31]) );
  DFFR_X1 out_reg_30_ ( .D(in[30]), .CK(clk), .RN(n2), .Q(out[30]) );
  DFFR_X1 out_reg_29_ ( .D(in[29]), .CK(clk), .RN(n2), .Q(out[29]) );
  DFFR_X1 out_reg_28_ ( .D(in[28]), .CK(clk), .RN(n2), .Q(out[28]) );
  DFFR_X1 out_reg_27_ ( .D(in[27]), .CK(clk), .RN(n2), .Q(out[27]) );
  DFFR_X1 out_reg_26_ ( .D(in[26]), .CK(clk), .RN(n2), .Q(out[26]) );
  DFFR_X1 out_reg_25_ ( .D(in[25]), .CK(clk), .RN(n2), .Q(out[25]) );
  DFFR_X1 out_reg_24_ ( .D(in[24]), .CK(clk), .RN(n2), .Q(out[24]) );
  DFFR_X1 out_reg_23_ ( .D(in[23]), .CK(clk), .RN(n2), .Q(out[23]) );
  DFFR_X1 out_reg_22_ ( .D(in[22]), .CK(clk), .RN(n2), .Q(out[22]) );
  DFFR_X1 out_reg_21_ ( .D(in[21]), .CK(clk), .RN(n2), .Q(out[21]) );
  DFFR_X1 out_reg_20_ ( .D(in[20]), .CK(clk), .RN(n2), .Q(out[20]) );
  DFFR_X1 out_reg_19_ ( .D(in[19]), .CK(clk), .RN(n2), .Q(out[19]) );
  DFFR_X1 out_reg_18_ ( .D(in[18]), .CK(clk), .RN(n2), .Q(out[18]) );
  DFFR_X1 out_reg_17_ ( .D(in[17]), .CK(clk), .RN(n2), .Q(out[17]) );
  DFFR_X1 out_reg_16_ ( .D(in[16]), .CK(clk), .RN(n2), .Q(out[16]) );
  DFFR_X1 out_reg_15_ ( .D(in[15]), .CK(clk), .RN(n2), .Q(out[15]) );
  DFFR_X1 out_reg_14_ ( .D(in[14]), .CK(clk), .RN(n2), .Q(out[14]) );
  DFFR_X1 out_reg_13_ ( .D(in[13]), .CK(clk), .RN(n2), .Q(out[13]) );
  DFFR_X1 out_reg_12_ ( .D(in[12]), .CK(clk), .RN(n2), .Q(out[12]) );
  DFFR_X1 out_reg_11_ ( .D(in[11]), .CK(clk), .RN(n2), .Q(out[11]) );
  DFFR_X1 out_reg_10_ ( .D(in[10]), .CK(clk), .RN(n2), .Q(out[10]) );
  DFFR_X1 out_reg_9_ ( .D(in[9]), .CK(clk), .RN(n2), .Q(out[9]) );
  DFFR_X1 out_reg_8_ ( .D(in[8]), .CK(clk), .RN(n2), .Q(out[8]) );
  DFFR_X1 out_reg_7_ ( .D(in[7]), .CK(clk), .RN(n2), .Q(out[7]) );
  DFFR_X1 out_reg_6_ ( .D(in[6]), .CK(clk), .RN(n2), .Q(out[6]) );
  DFFR_X1 out_reg_5_ ( .D(in[5]), .CK(clk), .RN(n2), .Q(out[5]) );
  DFFR_X1 out_reg_4_ ( .D(in[4]), .CK(clk), .RN(n2), .Q(out[4]) );
  DFFR_X1 out_reg_3_ ( .D(in[3]), .CK(clk), .RN(n2), .Q(out[3]) );
  DFFR_X1 out_reg_2_ ( .D(in[2]), .CK(clk), .RN(n2), .Q(out[2]) );
  DFFR_X1 out_reg_1_ ( .D(in[1]), .CK(clk), .RN(n2), .Q(out[1]) );
  DFFR_X1 out_reg_0_ ( .D(in[0]), .CK(clk), .RN(n2), .Q(out[0]) );
  INV_X4 U3 ( .A(rst), .ZN(n2) );
endmodule


module MUX2X1_0 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n3, n1;

  INV_X1 U1 ( .A(n3), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n3) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_114 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_113 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_112 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_111 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_110 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_109 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_108 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_107 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_106 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_105 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_104 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_103 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_102 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_101 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_100 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_99 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_98 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_97 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_96 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_95 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_94 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_93 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_92 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_91 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_90 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_89 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_88 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_87 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_86 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_85 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_84 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_83 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_82 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_81 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_80 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_79 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_78 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_77 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_76 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_75 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_74 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_73 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_72 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_71 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_70 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_69 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_68 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_67 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_66 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_65 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_64 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_63 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_62 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_61 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(n1), .A2(in0), .B1(in1), .B2(sel), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_60 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_59 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_58 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_57 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_56 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_55 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_54 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_53 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_52 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_51 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_50 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_49 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_48 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_47 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_46 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_45 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_44 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_43 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_42 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(in1), .B2(sel), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_41 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_40 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_39 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_38 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_37 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_36 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_35 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_34 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_33 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_32 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_31 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_30 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_29 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_28 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_27 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_26 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_25 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_24 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_23 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(out) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_22 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_21 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_20 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_19 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_18 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_17 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_16 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_15 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_14 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_13 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_12 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_11 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_10 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_9 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_8 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_7 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_6 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_5 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_4 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_3 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_2 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module MUX2X1_1 ( in0, in1, sel, out );
  input in0, in1, sel;
  output out;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(out) );
  AOI22_X1 U2 ( .A1(in0), .A2(n1), .B1(sel), .B2(in1), .ZN(n4) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module BarrelShifter ( In, Out, Shift );
  input [22:0] In;
  output [22:0] Out;
  input [4:0] Shift;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [22:0] a;
  wire   [22:0] a1;
  wire   [22:0] a2;
  wire   [22:0] a3;

  MUX2X1_0 b2_0__M ( .in0(In[0]), .in1(In[1]), .sel(n10), .out(a[0]) );
  MUX2X1_114 b2_1__M ( .in0(In[1]), .in1(In[2]), .sel(n9), .out(a[1]) );
  MUX2X1_113 b2_2__M ( .in0(In[2]), .in1(In[3]), .sel(n9), .out(a[2]) );
  MUX2X1_112 b2_3__M ( .in0(In[3]), .in1(In[4]), .sel(n9), .out(a[3]) );
  MUX2X1_111 b2_4__M ( .in0(In[4]), .in1(In[5]), .sel(n9), .out(a[4]) );
  MUX2X1_110 b2_5__M ( .in0(In[5]), .in1(In[6]), .sel(n9), .out(a[5]) );
  MUX2X1_109 b2_6__M ( .in0(In[6]), .in1(In[7]), .sel(n9), .out(a[6]) );
  MUX2X1_108 b2_7__M ( .in0(In[7]), .in1(In[8]), .sel(n9), .out(a[7]) );
  MUX2X1_107 b2_8__M ( .in0(In[8]), .in1(In[9]), .sel(n9), .out(a[8]) );
  MUX2X1_106 b2_9__M ( .in0(In[9]), .in1(In[10]), .sel(n9), .out(a[9]) );
  MUX2X1_105 b2_10__M ( .in0(In[10]), .in1(In[11]), .sel(n9), .out(a[10]) );
  MUX2X1_104 b2_11__M ( .in0(In[11]), .in1(In[12]), .sel(n9), .out(a[11]) );
  MUX2X1_103 b2_12__M ( .in0(In[12]), .in1(In[13]), .sel(n9), .out(a[12]) );
  MUX2X1_102 b2_13__M ( .in0(In[13]), .in1(In[14]), .sel(n10), .out(a[13]) );
  MUX2X1_101 b2_14__M ( .in0(In[14]), .in1(In[15]), .sel(n10), .out(a[14]) );
  MUX2X1_100 b2_15__M ( .in0(In[15]), .in1(In[16]), .sel(n10), .out(a[15]) );
  MUX2X1_99 b2_16__M ( .in0(In[16]), .in1(In[17]), .sel(n10), .out(a[16]) );
  MUX2X1_98 b2_17__M ( .in0(In[17]), .in1(In[18]), .sel(n10), .out(a[17]) );
  MUX2X1_97 b2_18__M ( .in0(In[18]), .in1(In[19]), .sel(n10), .out(a[18]) );
  MUX2X1_96 b2_19__M ( .in0(In[19]), .in1(In[20]), .sel(n10), .out(a[19]) );
  MUX2X1_95 b2_20__M ( .in0(In[20]), .in1(In[21]), .sel(n10), .out(a[20]) );
  MUX2X1_94 b2_21__M ( .in0(In[21]), .in1(In[22]), .sel(n10), .out(a[21]) );
  MUX2X1_93 M1 ( .in0(In[22]), .in1(1'b0), .sel(n10), .out(a[22]) );
  MUX2X1_92 b4_0__M2 ( .in0(a[0]), .in1(a[2]), .sel(n11), .out(a1[0]) );
  MUX2X1_91 b4_1__M2 ( .in0(a[1]), .in1(a[3]), .sel(n11), .out(a1[1]) );
  MUX2X1_90 b4_2__M2 ( .in0(a[2]), .in1(a[4]), .sel(n11), .out(a1[2]) );
  MUX2X1_89 b4_3__M2 ( .in0(a[3]), .in1(a[5]), .sel(n11), .out(a1[3]) );
  MUX2X1_88 b4_4__M2 ( .in0(a[4]), .in1(a[6]), .sel(n11), .out(a1[4]) );
  MUX2X1_87 b4_5__M2 ( .in0(a[5]), .in1(a[7]), .sel(n11), .out(a1[5]) );
  MUX2X1_86 b4_6__M2 ( .in0(a[6]), .in1(a[8]), .sel(n11), .out(a1[6]) );
  MUX2X1_85 b4_7__M2 ( .in0(a[7]), .in1(a[9]), .sel(n11), .out(a1[7]) );
  MUX2X1_84 b4_8__M2 ( .in0(a[8]), .in1(a[10]), .sel(n11), .out(a1[8]) );
  MUX2X1_83 b4_9__M2 ( .in0(a[9]), .in1(a[11]), .sel(n11), .out(a1[9]) );
  MUX2X1_82 b4_10__M2 ( .in0(a[10]), .in1(a[12]), .sel(n11), .out(a1[10]) );
  MUX2X1_81 b4_11__M2 ( .in0(a[11]), .in1(a[13]), .sel(n11), .out(a1[11]) );
  MUX2X1_80 b4_12__M2 ( .in0(a[12]), .in1(a[14]), .sel(n12), .out(a1[12]) );
  MUX2X1_79 b4_13__M2 ( .in0(a[13]), .in1(a[15]), .sel(n12), .out(a1[13]) );
  MUX2X1_78 b4_14__M2 ( .in0(a[14]), .in1(a[16]), .sel(n12), .out(a1[14]) );
  MUX2X1_77 b4_15__M2 ( .in0(a[15]), .in1(a[17]), .sel(n12), .out(a1[15]) );
  MUX2X1_76 b4_16__M2 ( .in0(a[16]), .in1(a[18]), .sel(n12), .out(a1[16]) );
  MUX2X1_75 b4_17__M2 ( .in0(a[17]), .in1(a[19]), .sel(n12), .out(a1[17]) );
  MUX2X1_74 b4_18__M2 ( .in0(a[18]), .in1(a[20]), .sel(n12), .out(a1[18]) );
  MUX2X1_73 b4_19__M2 ( .in0(a[19]), .in1(a[21]), .sel(n12), .out(a1[19]) );
  MUX2X1_72 b4_20__M2 ( .in0(a[20]), .in1(a[22]), .sel(n12), .out(a1[20]) );
  MUX2X1_71 b5_21__M3 ( .in0(a[21]), .in1(1'b0), .sel(n12), .out(a1[21]) );
  MUX2X1_70 b5_22__M3 ( .in0(a[22]), .in1(1'b0), .sel(n12), .out(a1[22]) );
  MUX2X1_69 b7_0__M4 ( .in0(a1[0]), .in1(a1[4]), .sel(n5), .out(a2[0]) );
  MUX2X1_68 b7_1__M4 ( .in0(a1[1]), .in1(a1[5]), .sel(n4), .out(a2[1]) );
  MUX2X1_67 b7_2__M4 ( .in0(a1[2]), .in1(a1[6]), .sel(n5), .out(a2[2]) );
  MUX2X1_66 b7_3__M4 ( .in0(a1[3]), .in1(a1[7]), .sel(n4), .out(a2[3]) );
  MUX2X1_65 b7_4__M4 ( .in0(a1[4]), .in1(a1[8]), .sel(n5), .out(a2[4]) );
  MUX2X1_64 b7_5__M4 ( .in0(a1[5]), .in1(a1[9]), .sel(n4), .out(a2[5]) );
  MUX2X1_63 b7_6__M4 ( .in0(a1[6]), .in1(a1[10]), .sel(n5), .out(a2[6]) );
  MUX2X1_62 b7_7__M4 ( .in0(a1[7]), .in1(a1[11]), .sel(n4), .out(a2[7]) );
  MUX2X1_61 b7_8__M4 ( .in0(a1[8]), .in1(a1[12]), .sel(n3), .out(a2[8]) );
  MUX2X1_60 b7_9__M4 ( .in0(a1[9]), .in1(a1[13]), .sel(n4), .out(a2[9]) );
  MUX2X1_59 b7_10__M4 ( .in0(a1[10]), .in1(a1[14]), .sel(n4), .out(a2[10]) );
  MUX2X1_58 b7_11__M4 ( .in0(a1[11]), .in1(a1[15]), .sel(n5), .out(a2[11]) );
  MUX2X1_57 b7_12__M4 ( .in0(a1[12]), .in1(a1[16]), .sel(n3), .out(a2[12]) );
  MUX2X1_56 b7_13__M4 ( .in0(a1[13]), .in1(a1[17]), .sel(n2), .out(a2[13]) );
  MUX2X1_55 b7_14__M4 ( .in0(a1[14]), .in1(a1[18]), .sel(n1), .out(a2[14]) );
  MUX2X1_54 b7_15__M4 ( .in0(a1[15]), .in1(a1[19]), .sel(n1), .out(a2[15]) );
  MUX2X1_53 b7_16__M4 ( .in0(a1[16]), .in1(a1[20]), .sel(n1), .out(a2[16]) );
  MUX2X1_52 b7_17__M4 ( .in0(a1[17]), .in1(a1[21]), .sel(n2), .out(a2[17]) );
  MUX2X1_51 b7_18__M4 ( .in0(a1[18]), .in1(a1[22]), .sel(n1), .out(a2[18]) );
  MUX2X1_50 b8_19__M5 ( .in0(a1[19]), .in1(1'b0), .sel(n2), .out(a2[19]) );
  MUX2X1_49 b8_20__M5 ( .in0(a1[20]), .in1(1'b0), .sel(n1), .out(a2[20]) );
  MUX2X1_48 b8_21__M5 ( .in0(a1[21]), .in1(1'b0), .sel(n2), .out(a2[21]) );
  MUX2X1_47 b8_22__M5 ( .in0(a1[22]), .in1(1'b0), .sel(n1), .out(a2[22]) );
  MUX2X1_46 b9_0__M6 ( .in0(a2[0]), .in1(a2[8]), .sel(n6), .out(a3[0]) );
  MUX2X1_45 b9_1__M6 ( .in0(a2[1]), .in1(a2[9]), .sel(n7), .out(a3[1]) );
  MUX2X1_44 b9_2__M6 ( .in0(a2[2]), .in1(a2[10]), .sel(n7), .out(a3[2]) );
  MUX2X1_43 b9_3__M6 ( .in0(a2[3]), .in1(a2[11]), .sel(n7), .out(a3[3]) );
  MUX2X1_42 b9_4__M6 ( .in0(a2[4]), .in1(a2[12]), .sel(n6), .out(a3[4]) );
  MUX2X1_41 b9_5__M6 ( .in0(a2[5]), .in1(a2[13]), .sel(n7), .out(a3[5]) );
  MUX2X1_40 b9_6__M6 ( .in0(a2[6]), .in1(a2[14]), .sel(n7), .out(a3[6]) );
  MUX2X1_39 b9_7__M6 ( .in0(a2[7]), .in1(a2[15]), .sel(n7), .out(a3[7]) );
  MUX2X1_38 b9_8__M6 ( .in0(a2[8]), .in1(a2[16]), .sel(n7), .out(a3[8]) );
  MUX2X1_37 b9_9__M6 ( .in0(a2[9]), .in1(a2[17]), .sel(n7), .out(a3[9]) );
  MUX2X1_36 b9_10__M6 ( .in0(a2[10]), .in1(a2[18]), .sel(n7), .out(a3[10]) );
  MUX2X1_35 b9_11__M6 ( .in0(a2[11]), .in1(a2[19]), .sel(n7), .out(a3[11]) );
  MUX2X1_34 b9_12__M6 ( .in0(a2[12]), .in1(a2[20]), .sel(n16), .out(a3[12]) );
  MUX2X1_33 b9_13__M6 ( .in0(a2[13]), .in1(a2[21]), .sel(n16), .out(a3[13]) );
  MUX2X1_32 b9_14__M6 ( .in0(a2[14]), .in1(a2[22]), .sel(n16), .out(a3[14]) );
  MUX2X1_31 b10_15__M7 ( .in0(a2[15]), .in1(1'b0), .sel(n16), .out(a3[15]) );
  MUX2X1_30 b10_16__M7 ( .in0(a2[16]), .in1(1'b0), .sel(n16), .out(a3[16]) );
  MUX2X1_29 b10_17__M7 ( .in0(a2[17]), .in1(1'b0), .sel(n16), .out(a3[17]) );
  MUX2X1_28 b10_18__M7 ( .in0(a2[18]), .in1(1'b0), .sel(n16), .out(a3[18]) );
  MUX2X1_27 b10_19__M7 ( .in0(a2[19]), .in1(1'b0), .sel(n16), .out(a3[19]) );
  MUX2X1_26 b10_20__M7 ( .in0(a2[20]), .in1(1'b0), .sel(n16), .out(a3[20]) );
  MUX2X1_25 b10_21__M7 ( .in0(a2[21]), .in1(1'b0), .sel(n16), .out(a3[21]) );
  MUX2X1_24 b10_22__M7 ( .in0(a2[22]), .in1(1'b0), .sel(n16), .out(a3[22]) );
  MUX2X1_23 b12_0__M8 ( .in0(a3[0]), .in1(a3[4]), .sel(Shift[4]), .out(Out[0])
         );
  MUX2X1_22 b12_1__M8 ( .in0(a3[1]), .in1(a3[5]), .sel(n8), .out(Out[1]) );
  MUX2X1_21 b12_2__M8 ( .in0(a3[2]), .in1(a3[6]), .sel(n8), .out(Out[2]) );
  MUX2X1_20 b12_3__M8 ( .in0(a3[3]), .in1(a3[7]), .sel(n8), .out(Out[3]) );
  MUX2X1_19 b12_4__M8 ( .in0(a3[4]), .in1(a3[8]), .sel(n8), .out(Out[4]) );
  MUX2X1_18 b12_5__M8 ( .in0(a3[5]), .in1(a3[9]), .sel(n8), .out(Out[5]) );
  MUX2X1_17 b12_6__M8 ( .in0(a3[6]), .in1(a3[10]), .sel(n8), .out(Out[6]) );
  MUX2X1_16 b13_7__M9 ( .in0(a3[7]), .in1(1'b0), .sel(n8), .out(Out[7]) );
  MUX2X1_15 b13_8__M9 ( .in0(a3[8]), .in1(1'b0), .sel(n8), .out(Out[8]) );
  MUX2X1_14 b13_9__M9 ( .in0(a3[9]), .in1(1'b0), .sel(n8), .out(Out[9]) );
  MUX2X1_13 b13_10__M9 ( .in0(a3[10]), .in1(1'b0), .sel(n8), .out(Out[10]) );
  MUX2X1_12 b13_11__M9 ( .in0(a3[11]), .in1(1'b0), .sel(n8), .out(Out[11]) );
  MUX2X1_11 b13_12__M9 ( .in0(a3[12]), .in1(1'b0), .sel(n18), .out(Out[12]) );
  MUX2X1_10 b13_13__M9 ( .in0(a3[13]), .in1(1'b0), .sel(n18), .out(Out[13]) );
  MUX2X1_9 b13_14__M9 ( .in0(a3[14]), .in1(1'b0), .sel(n18), .out(Out[14]) );
  MUX2X1_8 b13_15__M9 ( .in0(a3[15]), .in1(1'b0), .sel(n18), .out(Out[15]) );
  MUX2X1_7 b13_16__M9 ( .in0(a3[16]), .in1(1'b0), .sel(n18), .out(Out[16]) );
  MUX2X1_6 b13_17__M9 ( .in0(a3[17]), .in1(1'b0), .sel(n18), .out(Out[17]) );
  MUX2X1_5 b13_18__M9 ( .in0(a3[18]), .in1(1'b0), .sel(n18), .out(Out[18]) );
  MUX2X1_4 b13_19__M9 ( .in0(a3[19]), .in1(1'b0), .sel(n18), .out(Out[19]) );
  MUX2X1_3 b13_20__M9 ( .in0(a3[20]), .in1(1'b0), .sel(n18), .out(Out[20]) );
  MUX2X1_2 b13_21__M9 ( .in0(a3[21]), .in1(1'b0), .sel(n18), .out(Out[21]) );
  MUX2X1_1 b13_22__M9 ( .in0(a3[22]), .in1(1'b0), .sel(n18), .out(Out[22]) );
  BUF_X1 U2 ( .A(n13), .Z(n4) );
  BUF_X1 U3 ( .A(Shift[0]), .Z(n9) );
  BUF_X1 U4 ( .A(Shift[0]), .Z(n10) );
  CLKBUF_X3 U5 ( .A(n17), .Z(n8) );
  BUF_X2 U6 ( .A(n15), .Z(n7) );
  BUF_X1 U7 ( .A(n13), .Z(n5) );
  BUF_X1 U8 ( .A(n14), .Z(n2) );
  BUF_X1 U9 ( .A(n15), .Z(n6) );
  BUF_X2 U10 ( .A(Shift[1]), .Z(n11) );
  BUF_X2 U11 ( .A(Shift[1]), .Z(n12) );
  BUF_X1 U12 ( .A(Shift[2]), .Z(n13) );
  CLKBUF_X1 U13 ( .A(Shift[3]), .Z(n16) );
  BUF_X1 U14 ( .A(n14), .Z(n1) );
  BUF_X1 U15 ( .A(Shift[2]), .Z(n14) );
  CLKBUF_X1 U16 ( .A(n13), .Z(n3) );
  BUF_X1 U17 ( .A(Shift[3]), .Z(n15) );
  BUF_X1 U18 ( .A(Shift[4]), .Z(n17) );
  CLKBUF_X1 U19 ( .A(Shift[4]), .Z(n18) );
endmodule


module fpu_DW01_sub_23 ( A, B, CI, DIFF, CO );
  input [21:0] A;
  input [21:0] B;
  output [21:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;
  wire   [21:1] carry;

  FA_X1 U2_21 ( .A(A[21]), .B(n23), .CI(carry[21]), .S(DIFF[21]) );
  FA_X1 U2_20 ( .A(A[20]), .B(n22), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FA_X1 U2_19 ( .A(A[19]), .B(n21), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FA_X1 U2_18 ( .A(A[18]), .B(n20), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FA_X1 U2_17 ( .A(A[17]), .B(n19), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FA_X1 U2_16 ( .A(A[16]), .B(n18), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FA_X1 U2_15 ( .A(A[15]), .B(n17), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n16), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n15), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n14), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n13), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n12), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n11), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FA_X1 U2_8 ( .A(A[8]), .B(n10), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n9), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n8), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n7), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n4), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n3), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[1]), .ZN(n3) );
  NAND2_X1 U2 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U3 ( .A(A[0]), .ZN(n1) );
  INV_X1 U4 ( .A(B[2]), .ZN(n4) );
  INV_X1 U5 ( .A(B[3]), .ZN(n5) );
  INV_X1 U6 ( .A(B[4]), .ZN(n6) );
  INV_X1 U7 ( .A(B[5]), .ZN(n7) );
  INV_X1 U8 ( .A(B[6]), .ZN(n8) );
  XNOR2_X1 U9 ( .A(n2), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U10 ( .A(B[21]), .ZN(n23) );
  INV_X1 U11 ( .A(B[19]), .ZN(n21) );
  INV_X1 U12 ( .A(B[20]), .ZN(n22) );
  INV_X1 U13 ( .A(B[18]), .ZN(n20) );
  INV_X1 U14 ( .A(B[17]), .ZN(n19) );
  INV_X1 U15 ( .A(B[16]), .ZN(n18) );
  INV_X1 U16 ( .A(B[15]), .ZN(n17) );
  INV_X1 U17 ( .A(B[14]), .ZN(n16) );
  INV_X1 U18 ( .A(B[13]), .ZN(n15) );
  INV_X1 U19 ( .A(B[12]), .ZN(n14) );
  INV_X1 U20 ( .A(B[11]), .ZN(n13) );
  INV_X1 U21 ( .A(B[10]), .ZN(n12) );
  INV_X1 U22 ( .A(B[7]), .ZN(n9) );
  INV_X1 U23 ( .A(B[8]), .ZN(n10) );
  INV_X1 U24 ( .A(B[9]), .ZN(n11) );
  INV_X1 U25 ( .A(B[0]), .ZN(n2) );
endmodule


module fpu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [22:2] carry;

  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(SUM[23]), .S(SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module fpu ( in1, in2, overFlow, out );
  input [31:0] in1;
  input [31:0] in2;
  output [31:0] out;
  output overFlow;
  wire   N31, N97, N99, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N192, N193, N194, N195, N196, N197, N198,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N224, N225, N226, N229, N230, N231, N258, N259, N313, N314, N315,
         N316, N317, N318, N319, N320, N347, N348, N349, N350, N351, N352,
         N353, N354, N381, N382, N383, N384, N385, N386, N387, N388, N415,
         N416, N417, N418, N419, N420, N421, N422, N449, N450, N451, N452,
         N453, N454, N455, N456, N483, N484, N485, N486, N487, N488, N489,
         N490, N517, N518, N519, N520, N521, N522, N523, N524, N551, N552,
         N553, N554, N555, N556, N557, N558, N585, N586, N587, N588, N589,
         N590, N591, N592, N619, N620, N621, N622, N623, N624, N625, N626,
         N653, N654, N655, N656, N657, N658, N659, N660, N687, N688, N689,
         N690, N691, N692, N693, N694, N721, N722, N723, N724, N725, N726,
         N727, N728, N755, N756, N757, N758, N759, N760, N761, N762, N789,
         N790, N791, N792, N793, N794, N795, N796, N823, N824, N825, N826,
         N827, N828, N829, N830, N857, N858, N859, N860, N861, N862, N863,
         N864, N891, N892, N893, N894, N895, N896, N897, N898, N925, N926,
         N927, N928, N929, N930, N931, N932, N959, N960, N961, N962, N963,
         N964, N965, N966, N993, N994, N995, N996, N997, N998, N999, N1000,
         n3530, n3540, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n3810, n3820, n3830, n3840, n3850,
         n3860, n3870, n3880, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n4150, n4160, n4170, n4180,
         n4190, n4200, n4210, n4220, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n4490, n4500, n4510,
         n4520, n4530, n4540, n4550, n4560, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n4830, n4840,
         n4850, n4860, n4870, n4880, n4890, n4900, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n5170,
         n5180, n5190, n5200, n5210, n5220, n5230, n5240, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n5510, n5520, n5530, n5540, n5550, n5560, n5570, n5580, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n581, n582, n583,
         n584, n5850, n5860, n5870, n5880, n5890, n5900, n5910, n5920, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n6190, n6200, n6210, n6220, n6230, n6240, n6250,
         n6260, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n6530, n6540, n6550, n6560, n6570,
         n6580, n6590, n6600, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n6870, n6880, n6890, n6900,
         n6910, n6920, n6930, n6940, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n7210, n7220, n7230,
         n7240, n7250, n7260, n7270, n7280, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n7550, n7560,
         n7570, n7580, n7590, n7600, n7610, n7620, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n7890, n7900, n7910, n7920, n7930, n7940, n7950, n7960, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, sub_64_I22_aco_B_0_,
         sub_64_I21_aco_B_0_, sub_64_I20_aco_B_0_, sub_64_I19_aco_B_0_,
         sub_64_I18_aco_B_0_, sub_64_I17_aco_B_0_, sub_64_I16_aco_B_0_,
         sub_64_I15_aco_B_0_, sub_64_I14_aco_B_0_, sub_64_I13_aco_B_0_,
         sub_64_I12_aco_B_0_, sub_64_I11_aco_B_0_, sub_64_I10_aco_B_0_,
         sub_64_I9_aco_B_0_, sub_64_I8_aco_B_0_, sub_64_I7_aco_B_0_,
         sub_64_I6_aco_B_0_, sub_64_I5_aco_B_0_, sub_64_I4_aco_B_0_,
         sub_64_I3_aco_B_0_, sub_64_I2_aco_B_0_, sub_64_aco_B_0_,
         sub_64_aco_A_0_, sub_64_aco_A_1_, sub_64_aco_A_2_, sub_64_aco_A_5_,
         sub_64_aco_A_6_, sub_46_ni_B_0_, add_42_B_0_, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n3100, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n80, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n970, n98, n990, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n1740, n1750, n1760, n1770, n1780, n1790,
         n1800, n1810, n1820, n1830, n1840, n1850, n1860, n1870, n1880, n189,
         n190, n191, n1920, n1930, n1940, n1950, n1960, n1970, n1980, n199,
         n200, n2010, n2020, n2030, n2040, n2050, n2060, n2070, n2080, n2090,
         n2100, n2110, n2120, n2130, n2140, n2150, n2160, n2170, n2180, n2190,
         n2200, n2210, n2220, n223, n2240, n2250, n2260, n227, n228, n2290,
         n2300, n2310, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n2580, n2590, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n3101, n311, n312, n3130, n3140, n3150, n3160,
         n3170, n3180, n3190, n3200, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n3470, n3480, n3490,
         n3500, n3510, n3520, n355, n503, n541, n580, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n8230, n8240, n8250, n8260, n8270, n8280, n8290, n8300,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n8570, n8580, n8590, n8600, n8610, n8620,
         n8630, n8640, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n8910, n8920, n8930, n8940;
  wire   [30:0] a;
  wire   [27:0] b;
  wire   [4:0] shamt;
  wire   [22:0] inShift;
  wire   [7:0] Out_Exponent;
  wire   [7:1] sub_64_I22_aco_carry;
  wire   [7:1] sub_64_I21_aco_carry;
  wire   [7:1] sub_64_I20_aco_carry;
  wire   [7:1] sub_64_I19_aco_carry;
  wire   [7:1] sub_64_I18_aco_carry;
  wire   [7:1] sub_64_I17_aco_carry;
  wire   [7:1] sub_64_I16_aco_carry;
  wire   [7:1] sub_64_I15_aco_carry;
  wire   [7:1] sub_64_I14_aco_carry;
  wire   [7:1] sub_64_I13_aco_carry;
  wire   [7:1] sub_64_I12_aco_carry;
  wire   [7:1] sub_64_I11_aco_carry;
  wire   [7:1] sub_64_I10_aco_carry;
  wire   [7:1] sub_64_I9_aco_carry;
  wire   [7:1] sub_64_I8_aco_carry;
  wire   [7:1] sub_64_I7_aco_carry;
  wire   [7:1] sub_64_I6_aco_carry;
  wire   [7:1] sub_64_I5_aco_carry;
  wire   [7:1] sub_64_I4_aco_carry;
  wire   [7:1] sub_64_I3_aco_carry;
  wire   [7:1] sub_64_I2_aco_carry;
  wire   [7:1] sub_64_aco_carry;
  wire   [7:1] sub_46_ni_carry;
  wire   [7:2] add_42_carry;
  wire   [4:1] sub_36_carry;

  OAI21_X2 U569 ( .B1(n7960), .B2(n797), .A(n7910), .ZN(n630) );
  XOR2_X1 U857 ( .A(n66), .B(sub_64_I17_aco_B_0_), .Z(n507) );
  XOR2_X1 U858 ( .A(n78), .B(sub_64_I15_aco_B_0_), .Z(n5240) );
  XOR2_X1 U859 ( .A(n4550), .B(n582), .Z(n581) );
  XOR2_X1 U860 ( .A(n82), .B(n19), .Z(n548) );
  XOR2_X1 U861 ( .A(n80), .B(sub_64_I19_aco_B_0_), .Z(n4860) );
  BarrelShifter bs ( .In(inShift), .Out(b[22:0]), .Shift(shamt) );
  fpu_DW01_sub_23 sub_45 ( .A(a[21:0]), .B(b[21:0]), .CI(1'b0), .DIFF({N222, 
        N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, 
        N209, N208, N207, N206, N205, N204, N203, N202, N201}) );
  fpu_DW01_add_1 add_39 ( .A({1'b0, a[22:0]}), .B({1'b0, b[22:0]}), .CI(1'b0), 
        .SUM({N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, 
        N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, 
        N165}) );
  FA_X1 sub_36_U2_1 ( .A(a[24]), .B(n148), .CI(sub_36_carry[1]), .CO(
        sub_36_carry[2]), .S(shamt[1]) );
  FA_X1 sub_36_U2_2 ( .A(a[25]), .B(n149), .CI(sub_36_carry[2]), .CO(
        sub_36_carry[3]), .S(shamt[2]) );
  FA_X1 sub_36_U2_3 ( .A(a[26]), .B(n150), .CI(sub_36_carry[3]), .CO(
        sub_36_carry[4]), .S(shamt[3]) );
  FA_X1 sub_36_U2_4 ( .A(a[27]), .B(n151), .CI(sub_36_carry[4]), .S(shamt[4])
         );
  FA_X1 add_42_U1_7 ( .A(a[30]), .B(1'b0), .CI(add_42_carry[7]), .CO(overFlow), 
        .S(N198) );
  FA_X1 add_42_U1_6 ( .A(a[29]), .B(1'b0), .CI(add_42_carry[6]), .CO(
        add_42_carry[7]), .S(N197) );
  FA_X1 add_42_U1_5 ( .A(a[28]), .B(1'b0), .CI(add_42_carry[5]), .CO(
        add_42_carry[6]), .S(N196) );
  FA_X1 add_42_U1_4 ( .A(a[27]), .B(1'b0), .CI(add_42_carry[4]), .CO(
        add_42_carry[5]), .S(N195) );
  FA_X1 add_42_U1_3 ( .A(a[26]), .B(1'b0), .CI(add_42_carry[3]), .CO(
        add_42_carry[4]), .S(N194) );
  FA_X1 add_42_U1_2 ( .A(a[25]), .B(1'b0), .CI(add_42_carry[2]), .CO(
        add_42_carry[3]), .S(N193) );
  FA_X1 add_42_U1_1 ( .A(a[24]), .B(1'b0), .CI(n10), .CO(add_42_carry[2]), .S(
        N192) );
  FA_X1 sub_64_aco_U2_2 ( .A(sub_64_aco_A_2_), .B(1'b1), .CI(
        sub_64_aco_carry[2]), .CO(sub_64_aco_carry[3]), .S(N315) );
  FA_X1 sub_64_aco_U2_3 ( .A(N258), .B(1'b1), .CI(sub_64_aco_carry[3]), .CO(
        sub_64_aco_carry[4]), .S(N316) );
  FA_X1 sub_64_aco_U2_4 ( .A(N259), .B(1'b1), .CI(sub_64_aco_carry[4]), .CO(
        sub_64_aco_carry[5]), .S(N317) );
  FA_X1 sub_64_aco_U2_5 ( .A(sub_64_aco_A_5_), .B(1'b1), .CI(
        sub_64_aco_carry[5]), .CO(sub_64_aco_carry[6]), .S(N318) );
  FA_X1 sub_64_aco_U2_6 ( .A(sub_64_aco_A_6_), .B(1'b1), .CI(
        sub_64_aco_carry[6]), .CO(sub_64_aco_carry[7]), .S(N319) );
  FA_X1 sub_64_I2_aco_U2_1 ( .A(N314), .B(1'b1), .CI(sub_64_I2_aco_carry[1]), 
        .CO(sub_64_I2_aco_carry[2]), .S(N348) );
  FA_X1 sub_64_I2_aco_U2_2 ( .A(N315), .B(1'b1), .CI(sub_64_I2_aco_carry[2]), 
        .CO(sub_64_I2_aco_carry[3]), .S(N349) );
  FA_X1 sub_64_I2_aco_U2_3 ( .A(N316), .B(1'b1), .CI(sub_64_I2_aco_carry[3]), 
        .CO(sub_64_I2_aco_carry[4]), .S(N350) );
  FA_X1 sub_64_I2_aco_U2_4 ( .A(N317), .B(1'b1), .CI(sub_64_I2_aco_carry[4]), 
        .CO(sub_64_I2_aco_carry[5]), .S(N351) );
  FA_X1 sub_64_I2_aco_U2_5 ( .A(N318), .B(1'b1), .CI(sub_64_I2_aco_carry[5]), 
        .CO(sub_64_I2_aco_carry[6]), .S(N352) );
  FA_X1 sub_64_I2_aco_U2_6 ( .A(N319), .B(1'b1), .CI(sub_64_I2_aco_carry[6]), 
        .CO(sub_64_I2_aco_carry[7]), .S(N353) );
  FA_X1 sub_64_I3_aco_U2_2 ( .A(N349), .B(1'b1), .CI(sub_64_I3_aco_carry[2]), 
        .CO(sub_64_I3_aco_carry[3]), .S(N383) );
  FA_X1 sub_64_I3_aco_U2_3 ( .A(N350), .B(1'b1), .CI(sub_64_I3_aco_carry[3]), 
        .CO(sub_64_I3_aco_carry[4]), .S(N384) );
  FA_X1 sub_64_I3_aco_U2_4 ( .A(N351), .B(1'b1), .CI(sub_64_I3_aco_carry[4]), 
        .CO(sub_64_I3_aco_carry[5]), .S(N385) );
  FA_X1 sub_64_I3_aco_U2_5 ( .A(N352), .B(1'b1), .CI(sub_64_I3_aco_carry[5]), 
        .CO(sub_64_I3_aco_carry[6]), .S(N386) );
  FA_X1 sub_64_I3_aco_U2_6 ( .A(N353), .B(1'b1), .CI(sub_64_I3_aco_carry[6]), 
        .CO(sub_64_I3_aco_carry[7]), .S(N387) );
  FA_X1 sub_64_I4_aco_U2_1 ( .A(N382), .B(1'b1), .CI(sub_64_I4_aco_carry[1]), 
        .CO(sub_64_I4_aco_carry[2]), .S(N416) );
  FA_X1 sub_64_I4_aco_U2_2 ( .A(N383), .B(1'b1), .CI(sub_64_I4_aco_carry[2]), 
        .CO(sub_64_I4_aco_carry[3]), .S(N417) );
  FA_X1 sub_64_I4_aco_U2_3 ( .A(N384), .B(1'b1), .CI(sub_64_I4_aco_carry[3]), 
        .CO(sub_64_I4_aco_carry[4]), .S(N418) );
  FA_X1 sub_64_I4_aco_U2_4 ( .A(N385), .B(1'b1), .CI(sub_64_I4_aco_carry[4]), 
        .CO(sub_64_I4_aco_carry[5]), .S(N419) );
  FA_X1 sub_64_I4_aco_U2_5 ( .A(N386), .B(1'b1), .CI(sub_64_I4_aco_carry[5]), 
        .CO(sub_64_I4_aco_carry[6]), .S(N420) );
  FA_X1 sub_64_I4_aco_U2_6 ( .A(N387), .B(1'b1), .CI(sub_64_I4_aco_carry[6]), 
        .CO(sub_64_I4_aco_carry[7]), .S(N421) );
  FA_X1 sub_64_I5_aco_U2_2 ( .A(N417), .B(1'b1), .CI(sub_64_I5_aco_carry[2]), 
        .CO(sub_64_I5_aco_carry[3]), .S(N451) );
  FA_X1 sub_64_I5_aco_U2_3 ( .A(N418), .B(1'b1), .CI(sub_64_I5_aco_carry[3]), 
        .CO(sub_64_I5_aco_carry[4]), .S(N452) );
  FA_X1 sub_64_I5_aco_U2_4 ( .A(N419), .B(1'b1), .CI(sub_64_I5_aco_carry[4]), 
        .CO(sub_64_I5_aco_carry[5]), .S(N453) );
  FA_X1 sub_64_I5_aco_U2_5 ( .A(N420), .B(1'b1), .CI(sub_64_I5_aco_carry[5]), 
        .CO(sub_64_I5_aco_carry[6]), .S(N454) );
  FA_X1 sub_64_I5_aco_U2_6 ( .A(N421), .B(1'b1), .CI(sub_64_I5_aco_carry[6]), 
        .CO(sub_64_I5_aco_carry[7]), .S(N455) );
  FA_X1 sub_64_I6_aco_U2_1 ( .A(N450), .B(1'b1), .CI(sub_64_I6_aco_carry[1]), 
        .CO(sub_64_I6_aco_carry[2]), .S(N484) );
  FA_X1 sub_64_I6_aco_U2_2 ( .A(N451), .B(1'b1), .CI(sub_64_I6_aco_carry[2]), 
        .CO(sub_64_I6_aco_carry[3]), .S(N485) );
  FA_X1 sub_64_I6_aco_U2_3 ( .A(N452), .B(1'b1), .CI(sub_64_I6_aco_carry[3]), 
        .CO(sub_64_I6_aco_carry[4]), .S(N486) );
  FA_X1 sub_64_I6_aco_U2_4 ( .A(N453), .B(1'b1), .CI(sub_64_I6_aco_carry[4]), 
        .CO(sub_64_I6_aco_carry[5]), .S(N487) );
  FA_X1 sub_64_I6_aco_U2_5 ( .A(N454), .B(1'b1), .CI(sub_64_I6_aco_carry[5]), 
        .CO(sub_64_I6_aco_carry[6]), .S(N488) );
  FA_X1 sub_64_I6_aco_U2_6 ( .A(N455), .B(1'b1), .CI(sub_64_I6_aco_carry[6]), 
        .CO(sub_64_I6_aco_carry[7]), .S(N489) );
  FA_X1 sub_64_I7_aco_U2_2 ( .A(N485), .B(1'b1), .CI(sub_64_I7_aco_carry[2]), 
        .CO(sub_64_I7_aco_carry[3]), .S(N519) );
  FA_X1 sub_64_I7_aco_U2_3 ( .A(N486), .B(1'b1), .CI(sub_64_I7_aco_carry[3]), 
        .CO(sub_64_I7_aco_carry[4]), .S(N520) );
  FA_X1 sub_64_I7_aco_U2_4 ( .A(N487), .B(1'b1), .CI(sub_64_I7_aco_carry[4]), 
        .CO(sub_64_I7_aco_carry[5]), .S(N521) );
  FA_X1 sub_64_I7_aco_U2_5 ( .A(N488), .B(1'b1), .CI(sub_64_I7_aco_carry[5]), 
        .CO(sub_64_I7_aco_carry[6]), .S(N522) );
  FA_X1 sub_64_I7_aco_U2_6 ( .A(N489), .B(1'b1), .CI(sub_64_I7_aco_carry[6]), 
        .CO(sub_64_I7_aco_carry[7]), .S(N523) );
  FA_X1 sub_64_I8_aco_U2_1 ( .A(N518), .B(1'b1), .CI(sub_64_I8_aco_carry[1]), 
        .CO(sub_64_I8_aco_carry[2]), .S(N552) );
  FA_X1 sub_64_I8_aco_U2_2 ( .A(N519), .B(1'b1), .CI(sub_64_I8_aco_carry[2]), 
        .CO(sub_64_I8_aco_carry[3]), .S(N553) );
  FA_X1 sub_64_I8_aco_U2_3 ( .A(N520), .B(1'b1), .CI(sub_64_I8_aco_carry[3]), 
        .CO(sub_64_I8_aco_carry[4]), .S(N554) );
  FA_X1 sub_64_I8_aco_U2_4 ( .A(N521), .B(1'b1), .CI(sub_64_I8_aco_carry[4]), 
        .CO(sub_64_I8_aco_carry[5]), .S(N555) );
  FA_X1 sub_64_I8_aco_U2_5 ( .A(N522), .B(1'b1), .CI(sub_64_I8_aco_carry[5]), 
        .CO(sub_64_I8_aco_carry[6]), .S(N556) );
  FA_X1 sub_64_I8_aco_U2_6 ( .A(N523), .B(1'b1), .CI(sub_64_I8_aco_carry[6]), 
        .CO(sub_64_I8_aco_carry[7]), .S(N557) );
  FA_X1 sub_64_I9_aco_U2_2 ( .A(N553), .B(1'b1), .CI(sub_64_I9_aco_carry[2]), 
        .CO(sub_64_I9_aco_carry[3]), .S(N587) );
  FA_X1 sub_64_I9_aco_U2_3 ( .A(N554), .B(1'b1), .CI(sub_64_I9_aco_carry[3]), 
        .CO(sub_64_I9_aco_carry[4]), .S(N588) );
  FA_X1 sub_64_I9_aco_U2_4 ( .A(N555), .B(1'b1), .CI(sub_64_I9_aco_carry[4]), 
        .CO(sub_64_I9_aco_carry[5]), .S(N589) );
  FA_X1 sub_64_I9_aco_U2_5 ( .A(N556), .B(1'b1), .CI(sub_64_I9_aco_carry[5]), 
        .CO(sub_64_I9_aco_carry[6]), .S(N590) );
  FA_X1 sub_64_I9_aco_U2_6 ( .A(N557), .B(1'b1), .CI(sub_64_I9_aco_carry[6]), 
        .CO(sub_64_I9_aco_carry[7]), .S(N591) );
  FA_X1 sub_64_I10_aco_U2_1 ( .A(N586), .B(1'b1), .CI(sub_64_I10_aco_carry[1]), 
        .CO(sub_64_I10_aco_carry[2]), .S(N620) );
  FA_X1 sub_64_I10_aco_U2_2 ( .A(N587), .B(1'b1), .CI(sub_64_I10_aco_carry[2]), 
        .CO(sub_64_I10_aco_carry[3]), .S(N621) );
  FA_X1 sub_64_I10_aco_U2_3 ( .A(N588), .B(1'b1), .CI(sub_64_I10_aco_carry[3]), 
        .CO(sub_64_I10_aco_carry[4]), .S(N622) );
  FA_X1 sub_64_I10_aco_U2_4 ( .A(N589), .B(1'b1), .CI(sub_64_I10_aco_carry[4]), 
        .CO(sub_64_I10_aco_carry[5]), .S(N623) );
  FA_X1 sub_64_I10_aco_U2_5 ( .A(N590), .B(1'b1), .CI(sub_64_I10_aco_carry[5]), 
        .CO(sub_64_I10_aco_carry[6]), .S(N624) );
  FA_X1 sub_64_I10_aco_U2_6 ( .A(N591), .B(1'b1), .CI(sub_64_I10_aco_carry[6]), 
        .CO(sub_64_I10_aco_carry[7]), .S(N625) );
  FA_X1 sub_64_I11_aco_U2_2 ( .A(N621), .B(1'b1), .CI(sub_64_I11_aco_carry[2]), 
        .CO(sub_64_I11_aco_carry[3]), .S(N655) );
  FA_X1 sub_64_I11_aco_U2_3 ( .A(N622), .B(1'b1), .CI(sub_64_I11_aco_carry[3]), 
        .CO(sub_64_I11_aco_carry[4]), .S(N656) );
  FA_X1 sub_64_I11_aco_U2_4 ( .A(N623), .B(1'b1), .CI(sub_64_I11_aco_carry[4]), 
        .CO(sub_64_I11_aco_carry[5]), .S(N657) );
  FA_X1 sub_64_I11_aco_U2_5 ( .A(N624), .B(1'b1), .CI(sub_64_I11_aco_carry[5]), 
        .CO(sub_64_I11_aco_carry[6]), .S(N658) );
  FA_X1 sub_64_I11_aco_U2_6 ( .A(N625), .B(1'b1), .CI(sub_64_I11_aco_carry[6]), 
        .CO(sub_64_I11_aco_carry[7]), .S(N659) );
  FA_X1 sub_64_I12_aco_U2_1 ( .A(N654), .B(1'b1), .CI(sub_64_I12_aco_carry[1]), 
        .CO(sub_64_I12_aco_carry[2]), .S(N688) );
  FA_X1 sub_64_I12_aco_U2_2 ( .A(N655), .B(1'b1), .CI(sub_64_I12_aco_carry[2]), 
        .CO(sub_64_I12_aco_carry[3]), .S(N689) );
  FA_X1 sub_64_I12_aco_U2_3 ( .A(N656), .B(1'b1), .CI(sub_64_I12_aco_carry[3]), 
        .CO(sub_64_I12_aco_carry[4]), .S(N690) );
  FA_X1 sub_64_I12_aco_U2_4 ( .A(N657), .B(1'b1), .CI(sub_64_I12_aco_carry[4]), 
        .CO(sub_64_I12_aco_carry[5]), .S(N691) );
  FA_X1 sub_64_I12_aco_U2_5 ( .A(N658), .B(1'b1), .CI(sub_64_I12_aco_carry[5]), 
        .CO(sub_64_I12_aco_carry[6]), .S(N692) );
  FA_X1 sub_64_I12_aco_U2_6 ( .A(N659), .B(1'b1), .CI(sub_64_I12_aco_carry[6]), 
        .CO(sub_64_I12_aco_carry[7]), .S(N693) );
  FA_X1 sub_64_I13_aco_U2_2 ( .A(N689), .B(1'b1), .CI(sub_64_I13_aco_carry[2]), 
        .CO(sub_64_I13_aco_carry[3]), .S(N723) );
  FA_X1 sub_64_I13_aco_U2_3 ( .A(N690), .B(1'b1), .CI(sub_64_I13_aco_carry[3]), 
        .CO(sub_64_I13_aco_carry[4]), .S(N724) );
  FA_X1 sub_64_I13_aco_U2_4 ( .A(N691), .B(1'b1), .CI(sub_64_I13_aco_carry[4]), 
        .CO(sub_64_I13_aco_carry[5]), .S(N725) );
  FA_X1 sub_64_I13_aco_U2_5 ( .A(N692), .B(1'b1), .CI(sub_64_I13_aco_carry[5]), 
        .CO(sub_64_I13_aco_carry[6]), .S(N726) );
  FA_X1 sub_64_I13_aco_U2_6 ( .A(N693), .B(1'b1), .CI(sub_64_I13_aco_carry[6]), 
        .CO(sub_64_I13_aco_carry[7]), .S(N727) );
  FA_X1 sub_64_I14_aco_U2_1 ( .A(N722), .B(1'b1), .CI(sub_64_I14_aco_carry[1]), 
        .CO(sub_64_I14_aco_carry[2]), .S(N756) );
  FA_X1 sub_64_I14_aco_U2_2 ( .A(N723), .B(1'b1), .CI(sub_64_I14_aco_carry[2]), 
        .CO(sub_64_I14_aco_carry[3]), .S(N757) );
  FA_X1 sub_64_I14_aco_U2_3 ( .A(N724), .B(1'b1), .CI(sub_64_I14_aco_carry[3]), 
        .CO(sub_64_I14_aco_carry[4]), .S(N758) );
  FA_X1 sub_64_I14_aco_U2_4 ( .A(N725), .B(1'b1), .CI(sub_64_I14_aco_carry[4]), 
        .CO(sub_64_I14_aco_carry[5]), .S(N759) );
  FA_X1 sub_64_I14_aco_U2_5 ( .A(N726), .B(1'b1), .CI(sub_64_I14_aco_carry[5]), 
        .CO(sub_64_I14_aco_carry[6]), .S(N760) );
  FA_X1 sub_64_I14_aco_U2_6 ( .A(N727), .B(1'b1), .CI(sub_64_I14_aco_carry[6]), 
        .CO(sub_64_I14_aco_carry[7]), .S(N761) );
  FA_X1 sub_64_I15_aco_U2_2 ( .A(N757), .B(1'b1), .CI(sub_64_I15_aco_carry[2]), 
        .CO(sub_64_I15_aco_carry[3]), .S(N791) );
  FA_X1 sub_64_I15_aco_U2_3 ( .A(N758), .B(1'b1), .CI(sub_64_I15_aco_carry[3]), 
        .CO(sub_64_I15_aco_carry[4]), .S(N792) );
  FA_X1 sub_64_I15_aco_U2_4 ( .A(N759), .B(1'b1), .CI(sub_64_I15_aco_carry[4]), 
        .CO(sub_64_I15_aco_carry[5]), .S(N793) );
  FA_X1 sub_64_I15_aco_U2_5 ( .A(N760), .B(1'b1), .CI(sub_64_I15_aco_carry[5]), 
        .CO(sub_64_I15_aco_carry[6]), .S(N794) );
  FA_X1 sub_64_I15_aco_U2_6 ( .A(N761), .B(1'b1), .CI(sub_64_I15_aco_carry[6]), 
        .CO(sub_64_I15_aco_carry[7]), .S(N795) );
  FA_X1 sub_64_I16_aco_U2_1 ( .A(N790), .B(1'b1), .CI(sub_64_I16_aco_carry[1]), 
        .CO(sub_64_I16_aco_carry[2]), .S(N824) );
  FA_X1 sub_64_I16_aco_U2_2 ( .A(N791), .B(1'b1), .CI(sub_64_I16_aco_carry[2]), 
        .CO(sub_64_I16_aco_carry[3]), .S(N825) );
  FA_X1 sub_64_I16_aco_U2_3 ( .A(N792), .B(1'b1), .CI(sub_64_I16_aco_carry[3]), 
        .CO(sub_64_I16_aco_carry[4]), .S(N826) );
  FA_X1 sub_64_I16_aco_U2_4 ( .A(N793), .B(1'b1), .CI(sub_64_I16_aco_carry[4]), 
        .CO(sub_64_I16_aco_carry[5]), .S(N827) );
  FA_X1 sub_64_I16_aco_U2_5 ( .A(N794), .B(1'b1), .CI(sub_64_I16_aco_carry[5]), 
        .CO(sub_64_I16_aco_carry[6]), .S(N828) );
  FA_X1 sub_64_I16_aco_U2_6 ( .A(N795), .B(1'b1), .CI(sub_64_I16_aco_carry[6]), 
        .CO(sub_64_I16_aco_carry[7]), .S(N829) );
  FA_X1 sub_64_I17_aco_U2_2 ( .A(N825), .B(1'b1), .CI(sub_64_I17_aco_carry[2]), 
        .CO(sub_64_I17_aco_carry[3]), .S(N859) );
  FA_X1 sub_64_I17_aco_U2_3 ( .A(N826), .B(1'b1), .CI(sub_64_I17_aco_carry[3]), 
        .CO(sub_64_I17_aco_carry[4]), .S(N860) );
  FA_X1 sub_64_I17_aco_U2_4 ( .A(N827), .B(1'b1), .CI(sub_64_I17_aco_carry[4]), 
        .CO(sub_64_I17_aco_carry[5]), .S(N861) );
  FA_X1 sub_64_I17_aco_U2_5 ( .A(N828), .B(1'b1), .CI(sub_64_I17_aco_carry[5]), 
        .CO(sub_64_I17_aco_carry[6]), .S(N862) );
  FA_X1 sub_64_I17_aco_U2_6 ( .A(N829), .B(1'b1), .CI(sub_64_I17_aco_carry[6]), 
        .CO(sub_64_I17_aco_carry[7]), .S(N863) );
  FA_X1 sub_64_I18_aco_U2_1 ( .A(N858), .B(1'b1), .CI(sub_64_I18_aco_carry[1]), 
        .CO(sub_64_I18_aco_carry[2]), .S(N892) );
  FA_X1 sub_64_I18_aco_U2_2 ( .A(N859), .B(1'b1), .CI(sub_64_I18_aco_carry[2]), 
        .CO(sub_64_I18_aco_carry[3]), .S(N893) );
  FA_X1 sub_64_I18_aco_U2_3 ( .A(N860), .B(1'b1), .CI(sub_64_I18_aco_carry[3]), 
        .CO(sub_64_I18_aco_carry[4]), .S(N894) );
  FA_X1 sub_64_I18_aco_U2_4 ( .A(N861), .B(1'b1), .CI(sub_64_I18_aco_carry[4]), 
        .CO(sub_64_I18_aco_carry[5]), .S(N895) );
  FA_X1 sub_64_I18_aco_U2_5 ( .A(N862), .B(1'b1), .CI(sub_64_I18_aco_carry[5]), 
        .CO(sub_64_I18_aco_carry[6]), .S(N896) );
  FA_X1 sub_64_I18_aco_U2_6 ( .A(N863), .B(1'b1), .CI(sub_64_I18_aco_carry[6]), 
        .CO(sub_64_I18_aco_carry[7]), .S(N897) );
  FA_X1 sub_64_I19_aco_U2_1 ( .A(N892), .B(1'b1), .CI(sub_64_I19_aco_carry[1]), 
        .CO(sub_64_I19_aco_carry[2]), .S(N926) );
  FA_X1 sub_64_I19_aco_U2_2 ( .A(N893), .B(1'b1), .CI(sub_64_I19_aco_carry[2]), 
        .CO(sub_64_I19_aco_carry[3]), .S(N927) );
  FA_X1 sub_64_I19_aco_U2_3 ( .A(N894), .B(1'b1), .CI(sub_64_I19_aco_carry[3]), 
        .CO(sub_64_I19_aco_carry[4]), .S(N928) );
  FA_X1 sub_64_I19_aco_U2_4 ( .A(N895), .B(1'b1), .CI(sub_64_I19_aco_carry[4]), 
        .CO(sub_64_I19_aco_carry[5]), .S(N929) );
  FA_X1 sub_64_I19_aco_U2_5 ( .A(N896), .B(1'b1), .CI(sub_64_I19_aco_carry[5]), 
        .CO(sub_64_I19_aco_carry[6]), .S(N930) );
  FA_X1 sub_64_I19_aco_U2_6 ( .A(N897), .B(1'b1), .CI(sub_64_I19_aco_carry[6]), 
        .CO(sub_64_I19_aco_carry[7]), .S(N931) );
  FA_X1 sub_64_I20_aco_U2_1 ( .A(N926), .B(1'b1), .CI(sub_64_I20_aco_carry[1]), 
        .CO(sub_64_I20_aco_carry[2]), .S(N960) );
  FA_X1 sub_64_I20_aco_U2_2 ( .A(N927), .B(1'b1), .CI(sub_64_I20_aco_carry[2]), 
        .CO(sub_64_I20_aco_carry[3]), .S(N961) );
  FA_X1 sub_64_I20_aco_U2_3 ( .A(N928), .B(1'b1), .CI(sub_64_I20_aco_carry[3]), 
        .CO(sub_64_I20_aco_carry[4]), .S(N962) );
  FA_X1 sub_64_I20_aco_U2_4 ( .A(N929), .B(1'b1), .CI(sub_64_I20_aco_carry[4]), 
        .CO(sub_64_I20_aco_carry[5]), .S(N963) );
  FA_X1 sub_64_I20_aco_U2_5 ( .A(N930), .B(1'b1), .CI(sub_64_I20_aco_carry[5]), 
        .CO(sub_64_I20_aco_carry[6]), .S(N964) );
  FA_X1 sub_64_I20_aco_U2_6 ( .A(N931), .B(1'b1), .CI(sub_64_I20_aco_carry[6]), 
        .CO(sub_64_I20_aco_carry[7]), .S(N965) );
  FA_X1 sub_64_I21_aco_U2_2 ( .A(N961), .B(1'b1), .CI(sub_64_I21_aco_carry[2]), 
        .CO(sub_64_I21_aco_carry[3]), .S(N995) );
  FA_X1 sub_64_I21_aco_U2_3 ( .A(N962), .B(1'b1), .CI(sub_64_I21_aco_carry[3]), 
        .CO(sub_64_I21_aco_carry[4]), .S(N996) );
  FA_X1 sub_64_I21_aco_U2_4 ( .A(N963), .B(1'b1), .CI(sub_64_I21_aco_carry[4]), 
        .CO(sub_64_I21_aco_carry[5]), .S(N997) );
  FA_X1 sub_64_I21_aco_U2_5 ( .A(N964), .B(1'b1), .CI(sub_64_I21_aco_carry[5]), 
        .CO(sub_64_I21_aco_carry[6]), .S(N998) );
  FA_X1 sub_64_I21_aco_U2_6 ( .A(N965), .B(1'b1), .CI(sub_64_I21_aco_carry[6]), 
        .CO(sub_64_I21_aco_carry[7]), .S(N999) );
  FA_X1 sub_64_I22_aco_U2_1 ( .A(N994), .B(1'b1), .CI(sub_64_I22_aco_carry[1]), 
        .CO(sub_64_I22_aco_carry[2]), .S(Out_Exponent[1]) );
  FA_X1 sub_64_I22_aco_U2_2 ( .A(N995), .B(1'b1), .CI(sub_64_I22_aco_carry[2]), 
        .CO(sub_64_I22_aco_carry[3]), .S(Out_Exponent[2]) );
  FA_X1 sub_64_I22_aco_U2_3 ( .A(N996), .B(1'b1), .CI(sub_64_I22_aco_carry[3]), 
        .CO(sub_64_I22_aco_carry[4]), .S(Out_Exponent[3]) );
  FA_X1 sub_64_I22_aco_U2_4 ( .A(N997), .B(1'b1), .CI(sub_64_I22_aco_carry[4]), 
        .CO(sub_64_I22_aco_carry[5]), .S(Out_Exponent[4]) );
  FA_X1 sub_64_I22_aco_U2_5 ( .A(N998), .B(1'b1), .CI(sub_64_I22_aco_carry[5]), 
        .CO(sub_64_I22_aco_carry[6]), .S(Out_Exponent[5]) );
  FA_X1 sub_64_I22_aco_U2_6 ( .A(N999), .B(1'b1), .CI(sub_64_I22_aco_carry[6]), 
        .CO(sub_64_I22_aco_carry[7]), .S(Out_Exponent[6]) );
  AOI211_X1 U3 ( .C1(n841), .C2(n69), .A(n840), .B(n125), .ZN(n7910) );
  OAI221_X1 U4 ( .B1(n7940), .B2(n7950), .C1(n7900), .C2(n630), .A(n7910), 
        .ZN(n609) );
  OAI221_X1 U5 ( .B1(n7620), .B2(n763), .C1(n8290), .C2(n77), .A(n8300), .ZN(
        n571) );
  OAI21_X1 U6 ( .B1(n776), .B2(n777), .A(n768), .ZN(n6240) );
  OAI221_X1 U7 ( .B1(n749), .B2(n750), .C1(n737), .C2(n83), .A(n738), .ZN(
        n5520) );
  OAI221_X1 U8 ( .B1(n731), .B2(n732), .C1(n808), .C2(n76), .A(n809), .ZN(n530) );
  OAI221_X1 U9 ( .B1(n711), .B2(n712), .C1(n341), .C2(n82), .A(n342), .ZN(n511) );
  OAI221_X2 U10 ( .B1(n6880), .B2(n6890), .C1(n3180), .C2(n78), .A(n3190), 
        .ZN(n4900) );
  AOI22_X1 U11 ( .A1(N187), .A2(n129), .B1(N222), .B2(n136), .ZN(n370) );
  NAND2_X1 U12 ( .A1(n581), .A2(n837), .ZN(n469) );
  NAND2_X1 U13 ( .A1(n582), .A2(n837), .ZN(n3840) );
  BUF_X1 U14 ( .A(add_42_B_0_), .Z(n125) );
  XOR2_X2 U15 ( .A(n80), .B(n17), .Z(n389) );
  XOR2_X2 U16 ( .A(n66), .B(sub_64_I19_aco_B_0_), .Z(n395) );
  BUF_X1 U17 ( .A(n539), .Z(n105) );
  XOR2_X1 U18 ( .A(n603), .B(sub_64_I6_aco_B_0_), .Z(n1) );
  XOR2_X1 U19 ( .A(n628), .B(n606), .Z(n2) );
  BUF_X1 U20 ( .A(n85), .Z(n86) );
  NAND2_X1 U21 ( .A1(sub_64_I22_aco_B_0_), .A2(n837), .ZN(n3850) );
  XOR2_X1 U22 ( .A(n603), .B(sub_64_I6_aco_B_0_), .Z(n3) );
  XOR2_X1 U23 ( .A(n609), .B(sub_64_I2_aco_B_0_), .Z(n4) );
  XOR2_X1 U24 ( .A(n628), .B(n606), .Z(n5) );
  OR4_X1 U25 ( .A1(N997), .A2(N996), .A3(N999), .A4(N998), .ZN(n636) );
  OR4_X1 U26 ( .A1(N892), .A2(N891), .A3(N894), .A4(N893), .ZN(n666) );
  OR4_X1 U27 ( .A1(N348), .A2(N347), .A3(N350), .A4(N349), .ZN(n7950) );
  OR4_X1 U28 ( .A1(N416), .A2(N415), .A3(N418), .A4(N417), .ZN(n786) );
  OR4_X1 U29 ( .A1(N960), .A2(N959), .A3(N962), .A4(N961), .ZN(n640) );
  OR4_X1 U30 ( .A1(N688), .A2(N687), .A3(N690), .A4(N689), .ZN(n732) );
  OR4_X1 U31 ( .A1(N858), .A2(N857), .A3(N860), .A4(N859), .ZN(n668) );
  OR4_X1 U32 ( .A1(N824), .A2(N823), .A3(N826), .A4(N825), .ZN(n6890) );
  OR4_X1 U33 ( .A1(N484), .A2(N483), .A3(N486), .A4(N485), .ZN(n775) );
  OR4_X1 U34 ( .A1(N756), .A2(N755), .A3(N758), .A4(N757), .ZN(n712) );
  OR4_X1 U35 ( .A1(N620), .A2(N619), .A3(N622), .A4(N621), .ZN(n750) );
  OR4_X1 U36 ( .A1(N552), .A2(N551), .A3(N554), .A4(N553), .ZN(n763) );
  OR2_X1 U37 ( .A1(a[28]), .A2(sub_46_ni_carry[5]), .ZN(sub_46_ni_carry[6]) );
  XOR2_X1 U38 ( .A(n362), .B(n805), .Z(n6) );
  BUF_X1 U39 ( .A(n664), .Z(n88) );
  BUF_X1 U40 ( .A(n664), .Z(n87) );
  INV_X1 U41 ( .A(n445), .ZN(n275) );
  BUF_X1 U42 ( .A(n664), .Z(n89) );
  INV_X1 U43 ( .A(n6190), .ZN(n8270) );
  INV_X1 U44 ( .A(n643), .ZN(n274) );
  OAI221_X1 U45 ( .B1(n294), .B2(n394), .C1(n295), .C2(n395), .A(n296), .ZN(
        n643) );
  INV_X1 U46 ( .A(n715), .ZN(n342) );
  OAI221_X1 U47 ( .B1(n807), .B2(n424), .C1(n808), .C2(n425), .A(n809), .ZN(
        n715) );
  INV_X1 U49 ( .A(sub_64_aco_carry[1]), .ZN(n11) );
  NOR2_X1 U51 ( .A1(n70), .A2(n125), .ZN(n664) );
  OAI222_X1 U52 ( .A1(n300), .A2(n393), .B1(n3101), .B2(n394), .C1(n299), .C2(
        n395), .ZN(n445) );
  OAI22_X1 U53 ( .A1(n4860), .A2(n5870), .B1(n292), .B2(n4850), .ZN(n583) );
  INV_X1 U54 ( .A(n645), .ZN(n272) );
  OAI222_X1 U55 ( .A1(n294), .A2(n393), .B1(n297), .B2(n394), .C1(n298), .C2(
        n395), .ZN(n645) );
  INV_X1 U56 ( .A(n446), .ZN(n276) );
  OAI222_X1 U57 ( .A1(n301), .A2(n393), .B1(n299), .B2(n394), .C1(n300), .C2(
        n395), .ZN(n446) );
  INV_X1 U58 ( .A(n432), .ZN(n277) );
  OAI222_X1 U59 ( .A1(n302), .A2(n393), .B1(n300), .B2(n394), .C1(n301), .C2(
        n395), .ZN(n432) );
  INV_X1 U60 ( .A(n427), .ZN(n278) );
  OAI222_X1 U61 ( .A1(n303), .A2(n393), .B1(n301), .B2(n394), .C1(n302), .C2(
        n395), .ZN(n427) );
  INV_X1 U62 ( .A(n4190), .ZN(n279) );
  OAI222_X1 U63 ( .A1(n304), .A2(n393), .B1(n302), .B2(n394), .C1(n303), .C2(
        n395), .ZN(n4190) );
  INV_X1 U64 ( .A(n4150), .ZN(n280) );
  OAI222_X1 U65 ( .A1(n305), .A2(n393), .B1(n303), .B2(n394), .C1(n304), .C2(
        n395), .ZN(n4150) );
  INV_X1 U66 ( .A(n408), .ZN(n281) );
  OAI222_X1 U67 ( .A1(n306), .A2(n393), .B1(n304), .B2(n394), .C1(n305), .C2(
        n395), .ZN(n408) );
  INV_X1 U68 ( .A(n405), .ZN(n282) );
  OAI222_X1 U69 ( .A1(n307), .A2(n393), .B1(n305), .B2(n394), .C1(n306), .C2(
        n395), .ZN(n405) );
  INV_X1 U70 ( .A(n399), .ZN(n283) );
  OAI222_X1 U71 ( .A1(n308), .A2(n393), .B1(n306), .B2(n394), .C1(n307), .C2(
        n395), .ZN(n399) );
  INV_X1 U72 ( .A(n397), .ZN(n284) );
  OAI222_X1 U73 ( .A1(n297), .A2(n393), .B1(n307), .B2(n394), .C1(n308), .C2(
        n395), .ZN(n397) );
  INV_X1 U74 ( .A(n392), .ZN(n285) );
  OAI222_X1 U75 ( .A1(n298), .A2(n393), .B1(n308), .B2(n394), .C1(n297), .C2(
        n395), .ZN(n392) );
  INV_X1 U76 ( .A(n638), .ZN(n250) );
  OAI221_X1 U77 ( .B1(n272), .B2(n3880), .C1(n273), .C2(n389), .A(n274), .ZN(
        n638) );
  INV_X1 U78 ( .A(n4840), .ZN(n270) );
  OAI222_X1 U79 ( .A1(n287), .A2(n4850), .B1(n290), .B2(n471), .C1(n291), .C2(
        n4860), .ZN(n4840) );
  INV_X1 U80 ( .A(n5860), .ZN(n265) );
  OAI222_X1 U81 ( .A1(n293), .A2(n4850), .B1(n471), .B2(n5870), .C1(n292), 
        .C2(n4860), .ZN(n5860) );
  INV_X1 U82 ( .A(n5570), .ZN(n266) );
  OAI222_X1 U83 ( .A1(n288), .A2(n4850), .B1(n292), .B2(n471), .C1(n293), .C2(
        n4860), .ZN(n5570) );
  INV_X1 U84 ( .A(n542), .ZN(n267) );
  OAI222_X1 U85 ( .A1(n289), .A2(n4850), .B1(n293), .B2(n471), .C1(n288), .C2(
        n4860), .ZN(n542) );
  INV_X1 U86 ( .A(n5200), .ZN(n268) );
  OAI222_X1 U87 ( .A1(n290), .A2(n4850), .B1(n288), .B2(n471), .C1(n289), .C2(
        n4860), .ZN(n5200) );
  INV_X1 U88 ( .A(n504), .ZN(n269) );
  OAI222_X1 U89 ( .A1(n291), .A2(n4850), .B1(n289), .B2(n471), .C1(n290), .C2(
        n4860), .ZN(n504) );
  INV_X1 U90 ( .A(n644), .ZN(n273) );
  OAI222_X1 U91 ( .A1(n295), .A2(n393), .B1(n298), .B2(n394), .C1(n294), .C2(
        n395), .ZN(n644) );
  INV_X1 U92 ( .A(n6920), .ZN(n3190) );
  OAI221_X1 U93 ( .B1(n340), .B2(n412), .C1(n341), .C2(n413), .A(n342), .ZN(
        n6920) );
  INV_X1 U94 ( .A(n780), .ZN(n834) );
  INV_X1 U95 ( .A(n7550), .ZN(n8300) );
  INV_X1 U96 ( .A(n615), .ZN(n333) );
  INV_X1 U97 ( .A(n510), .ZN(n335) );
  AOI222_X1 U98 ( .A1(n125), .A2(n849), .B1(n851), .B2(n71), .C1(n850), .C2(
        n88), .ZN(n748) );
  AOI222_X1 U99 ( .A1(n125), .A2(n850), .B1(n852), .B2(n73), .C1(n851), .C2(
        n89), .ZN(n7280) );
  AOI222_X1 U100 ( .A1(n125), .A2(n851), .B1(n853), .B2(n74), .C1(n852), .C2(
        n88), .ZN(n729) );
  AOI222_X1 U101 ( .A1(n125), .A2(n852), .B1(n854), .B2(n75), .C1(n853), .C2(
        n87), .ZN(n707) );
  NAND2_X1 U102 ( .A1(n6220), .A2(n113), .ZN(n6190) );
  AOI222_X1 U103 ( .A1(n125), .A2(n8580), .B1(n8600), .B2(n71), .C1(n8590), 
        .C2(n88), .ZN(n575) );
  INV_X1 U104 ( .A(n577), .ZN(n835) );
  INV_X1 U105 ( .A(n631), .ZN(n836) );
  OAI222_X1 U106 ( .A1(n271), .A2(n4520), .B1(n265), .B2(n469), .C1(n266), 
        .C2(n470), .ZN(out[3]) );
  INV_X1 U107 ( .A(n583), .ZN(n271) );
  OAI222_X1 U108 ( .A1(n265), .A2(n4520), .B1(n266), .B2(n469), .C1(n267), 
        .C2(n470), .ZN(out[4]) );
  OAI222_X1 U109 ( .A1(n266), .A2(n4520), .B1(n267), .B2(n469), .C1(n268), 
        .C2(n470), .ZN(out[5]) );
  OAI222_X1 U110 ( .A1(n267), .A2(n4520), .B1(n268), .B2(n469), .C1(n269), 
        .C2(n470), .ZN(out[6]) );
  OAI222_X1 U111 ( .A1(n268), .A2(n4520), .B1(n269), .B2(n469), .C1(n270), 
        .C2(n470), .ZN(out[7]) );
  OAI222_X1 U112 ( .A1(n269), .A2(n4520), .B1(n270), .B2(n469), .C1(n264), 
        .C2(n470), .ZN(out[8]) );
  INV_X1 U113 ( .A(n4540), .ZN(n264) );
  INV_X1 U114 ( .A(n146), .ZN(n143) );
  OAI221_X1 U115 ( .B1(n265), .B2(n470), .C1(n584), .C2(n3850), .A(n5850), 
        .ZN(out[2]) );
  INV_X1 U116 ( .A(n3840), .ZN(n249) );
  OR2_X1 U117 ( .A1(n609), .A2(N347), .ZN(sub_64_I3_aco_carry[1]) );
  OR2_X1 U118 ( .A1(n4550), .A2(N959), .ZN(sub_64_I21_aco_carry[1]) );
  OR2_X1 U119 ( .A1(n634), .A2(sub_64_aco_A_0_), .ZN(sub_64_aco_carry[1]) );
  AOI222_X1 U120 ( .A1(n125), .A2(n841), .B1(n843), .B2(n73), .C1(n842), .C2(
        n87), .ZN(n7890) );
  AOI222_X1 U121 ( .A1(n125), .A2(n840), .B1(n842), .B2(n71), .C1(n841), .C2(
        n88), .ZN(n7900) );
  NAND2_X1 U122 ( .A1(sub_64_I11_aco_B_0_), .A2(sub_64_I10_aco_B_0_), .ZN(n440) );
  AOI222_X1 U123 ( .A1(n753), .A2(n114), .B1(n742), .B2(n466), .C1(n741), .C2(
        n468), .ZN(n736) );
  AOI222_X1 U124 ( .A1(n778), .A2(n96), .B1(n770), .B2(n104), .C1(n769), .C2(
        n2), .ZN(n766) );
  AOI222_X1 U125 ( .A1(n754), .A2(n115), .B1(n741), .B2(n466), .C1(n753), .C2(
        n468), .ZN(n737) );
  AOI222_X1 U126 ( .A1(n779), .A2(n970), .B1(n769), .B2(n106), .C1(n778), .C2(
        n5), .ZN(n767) );
  AOI221_X1 U127 ( .B1(n778), .B2(n105), .C1(n779), .C2(n2), .A(n780), .ZN(
        n768) );
  AOI221_X1 U128 ( .B1(n753), .B2(n466), .C1(n754), .C2(n468), .A(n7550), .ZN(
        n738) );
  OAI222_X1 U129 ( .A1(n7890), .A2(n90), .B1(n782), .B2(n91), .C1(n781), .C2(
        n86), .ZN(n778) );
  OAI222_X1 U130 ( .A1(n7900), .A2(n576), .B1(n781), .B2(n578), .C1(n7890), 
        .C2(n4), .ZN(n779) );
  OAI222_X1 U131 ( .A1(n766), .A2(n107), .B1(n7570), .B2(n108), .C1(n7560), 
        .C2(n1), .ZN(n753) );
  OAI222_X1 U132 ( .A1(n767), .A2(n499), .B1(n7560), .B2(n109), .C1(n766), 
        .C2(n3), .ZN(n754) );
  OAI221_X1 U133 ( .B1(n7890), .B2(n578), .C1(n7900), .C2(n86), .A(n7910), 
        .ZN(n780) );
  XNOR2_X1 U134 ( .A(n634), .B(sub_64_aco_A_0_), .ZN(N313) );
  OAI221_X1 U135 ( .B1(n766), .B2(n109), .C1(n767), .C2(n1), .A(n768), .ZN(
        n7550) );
  XNOR2_X1 U136 ( .A(n609), .B(N347), .ZN(N381) );
  XNOR2_X1 U137 ( .A(n66), .B(N857), .ZN(N891) );
  NAND2_X1 U138 ( .A1(n80), .A2(n15), .ZN(n4850) );
  XNOR2_X1 U139 ( .A(n4550), .B(N959), .ZN(N993) );
  NOR2_X1 U140 ( .A1(sub_64_I5_aco_B_0_), .A2(sub_64_I4_aco_B_0_), .ZN(n92) );
  INV_X1 U141 ( .A(n77), .ZN(sub_64_I8_aco_B_0_) );
  NOR2_X1 U142 ( .A1(n67), .A2(sub_64_I8_aco_B_0_), .ZN(n110) );
  NOR2_X1 U143 ( .A1(n3840), .A2(n611), .ZN(out[0]) );
  OAI22_X1 U144 ( .A1(n251), .A2(n3840), .B1(n443), .B2(n3850), .ZN(out[10])
         );
  OAI22_X1 U145 ( .A1(n252), .A2(n3840), .B1(n251), .B2(n3850), .ZN(out[11])
         );
  OAI22_X1 U146 ( .A1(n253), .A2(n3840), .B1(n252), .B2(n3850), .ZN(out[12])
         );
  OAI22_X1 U147 ( .A1(n254), .A2(n3840), .B1(n253), .B2(n3850), .ZN(out[13])
         );
  OAI22_X1 U148 ( .A1(n255), .A2(n3840), .B1(n254), .B2(n3850), .ZN(out[14])
         );
  OAI22_X1 U149 ( .A1(n256), .A2(n3840), .B1(n255), .B2(n3850), .ZN(out[15])
         );
  OAI22_X1 U150 ( .A1(n257), .A2(n3840), .B1(n256), .B2(n3850), .ZN(out[16])
         );
  OAI22_X1 U151 ( .A1(n2580), .A2(n3840), .B1(n257), .B2(n3850), .ZN(out[17])
         );
  OAI22_X1 U152 ( .A1(n2590), .A2(n3840), .B1(n2580), .B2(n3850), .ZN(out[18])
         );
  OAI22_X1 U153 ( .A1(n260), .A2(n3840), .B1(n2590), .B2(n3850), .ZN(out[19])
         );
  OAI22_X1 U154 ( .A1(n261), .A2(n3840), .B1(n260), .B2(n3850), .ZN(out[20])
         );
  OAI22_X1 U155 ( .A1(n262), .A2(n3840), .B1(n261), .B2(n3850), .ZN(out[21])
         );
  OAI22_X1 U156 ( .A1(n250), .A2(n3840), .B1(n262), .B2(n3850), .ZN(out[22])
         );
  OAI22_X1 U157 ( .A1(n584), .A2(n3840), .B1(n3850), .B2(n611), .ZN(out[1]) );
  INV_X1 U158 ( .A(n717), .ZN(n340) );
  OAI222_X1 U159 ( .A1(n807), .A2(n423), .B1(n810), .B2(n424), .C1(n811), .C2(
        n425), .ZN(n717) );
  BUF_X1 U160 ( .A(n539), .Z(n104) );
  INV_X1 U161 ( .A(n671), .ZN(n294) );
  OAI222_X1 U162 ( .A1(n3170), .A2(n401), .B1(n3200), .B2(n402), .C1(n321), 
        .C2(n403), .ZN(n671) );
  INV_X1 U163 ( .A(n6940), .ZN(n3170) );
  OAI222_X1 U164 ( .A1(n340), .A2(n411), .B1(n343), .B2(n412), .C1(n344), .C2(
        n413), .ZN(n6940) );
  INV_X1 U165 ( .A(n716), .ZN(n341) );
  OAI222_X1 U166 ( .A1(n808), .A2(n423), .B1(n811), .B2(n424), .C1(n807), .C2(
        n425), .ZN(n716) );
  INV_X1 U167 ( .A(n735), .ZN(n809) );
  OAI221_X1 U168 ( .B1(n736), .B2(n440), .C1(n737), .C2(n442), .A(n738), .ZN(
        n735) );
  INV_X1 U169 ( .A(n740), .ZN(n807) );
  OAI222_X1 U170 ( .A1(n736), .A2(n124), .B1(n720), .B2(n440), .C1(n719), .C2(
        n442), .ZN(n740) );
  INV_X1 U171 ( .A(n670), .ZN(n295) );
  OAI222_X1 U172 ( .A1(n3180), .A2(n401), .B1(n321), .B2(n402), .C1(n3170), 
        .C2(n403), .ZN(n670) );
  CLKBUF_X1 U173 ( .A(n539), .Z(n106) );
  INV_X1 U174 ( .A(n669), .ZN(n296) );
  OAI221_X1 U175 ( .B1(n3170), .B2(n402), .C1(n3180), .C2(n403), .A(n3190), 
        .ZN(n669) );
  INV_X1 U176 ( .A(n6930), .ZN(n3180) );
  OAI222_X1 U177 ( .A1(n341), .A2(n411), .B1(n344), .B2(n412), .C1(n340), .C2(
        n413), .ZN(n6930) );
  INV_X1 U178 ( .A(n739), .ZN(n808) );
  OAI222_X1 U179 ( .A1(n737), .A2(n124), .B1(n719), .B2(n440), .C1(n736), .C2(
        n442), .ZN(n739) );
  INV_X1 U180 ( .A(n376), .ZN(n841) );
  INV_X1 U181 ( .A(n444), .ZN(n251) );
  OAI222_X1 U182 ( .A1(n276), .A2(n3870), .B1(n286), .B2(n3880), .C1(n275), 
        .C2(n389), .ZN(n444) );
  INV_X1 U183 ( .A(n431), .ZN(n252) );
  OAI222_X1 U184 ( .A1(n277), .A2(n3870), .B1(n275), .B2(n3880), .C1(n276), 
        .C2(n389), .ZN(n431) );
  INV_X1 U185 ( .A(n426), .ZN(n253) );
  OAI222_X1 U186 ( .A1(n278), .A2(n3870), .B1(n276), .B2(n3880), .C1(n277), 
        .C2(n389), .ZN(n426) );
  INV_X1 U187 ( .A(n4180), .ZN(n254) );
  OAI222_X1 U188 ( .A1(n279), .A2(n3870), .B1(n277), .B2(n3880), .C1(n278), 
        .C2(n389), .ZN(n4180) );
  INV_X1 U189 ( .A(n414), .ZN(n255) );
  OAI222_X1 U190 ( .A1(n280), .A2(n3870), .B1(n278), .B2(n3880), .C1(n279), 
        .C2(n389), .ZN(n414) );
  INV_X1 U191 ( .A(n407), .ZN(n256) );
  OAI222_X1 U192 ( .A1(n281), .A2(n3870), .B1(n279), .B2(n3880), .C1(n280), 
        .C2(n389), .ZN(n407) );
  INV_X1 U193 ( .A(n404), .ZN(n257) );
  OAI222_X1 U194 ( .A1(n282), .A2(n3870), .B1(n280), .B2(n3880), .C1(n281), 
        .C2(n389), .ZN(n404) );
  INV_X1 U195 ( .A(n398), .ZN(n2580) );
  OAI222_X1 U196 ( .A1(n283), .A2(n3870), .B1(n281), .B2(n3880), .C1(n282), 
        .C2(n389), .ZN(n398) );
  INV_X1 U197 ( .A(n396), .ZN(n2590) );
  OAI222_X1 U198 ( .A1(n284), .A2(n3870), .B1(n282), .B2(n3880), .C1(n283), 
        .C2(n389), .ZN(n396) );
  INV_X1 U199 ( .A(n391), .ZN(n260) );
  OAI222_X1 U200 ( .A1(n285), .A2(n3870), .B1(n283), .B2(n3880), .C1(n284), 
        .C2(n389), .ZN(n391) );
  INV_X1 U201 ( .A(n390), .ZN(n261) );
  OAI222_X1 U202 ( .A1(n272), .A2(n3870), .B1(n284), .B2(n3880), .C1(n285), 
        .C2(n389), .ZN(n390) );
  INV_X1 U203 ( .A(n3860), .ZN(n262) );
  OAI222_X1 U204 ( .A1(n273), .A2(n3870), .B1(n285), .B2(n3880), .C1(n272), 
        .C2(n389), .ZN(n3860) );
  BUF_X1 U205 ( .A(n438), .Z(n124) );
  INV_X1 U206 ( .A(n3850), .ZN(n248) );
  XOR2_X1 U207 ( .A(add_42_B_0_), .B(n84), .Z(n7) );
  OAI221_X1 U208 ( .B1(n291), .B2(n471), .C1(sub_64_I20_aco_B_0_), .C2(n286), 
        .A(n472), .ZN(n4540) );
  AOI221_X1 U209 ( .B1(n445), .B2(n263), .C1(n4540), .C2(n17), .A(n4560), .ZN(
        n443) );
  INV_X1 U210 ( .A(n3870), .ZN(n263) );
  AOI222_X1 U211 ( .A1(n125), .A2(n842), .B1(n844), .B2(n74), .C1(n843), .C2(
        n89), .ZN(n781) );
  AOI222_X1 U212 ( .A1(n125), .A2(n843), .B1(n845), .B2(n75), .C1(n844), .C2(
        n89), .ZN(n782) );
  AOI222_X1 U213 ( .A1(n741), .A2(n119), .B1(n7220), .B2(n466), .C1(n742), 
        .C2(n468), .ZN(n719) );
  AOI222_X1 U214 ( .A1(n742), .A2(n118), .B1(n7230), .B2(n466), .C1(n7220), 
        .C2(n468), .ZN(n720) );
  AOI222_X1 U215 ( .A1(n769), .A2(n990), .B1(n7580), .B2(n105), .C1(n770), 
        .C2(n2), .ZN(n7560) );
  AOI222_X1 U216 ( .A1(n770), .A2(n98), .B1(n7590), .B2(n105), .C1(n7580), 
        .C2(n5), .ZN(n7570) );
  OAI222_X1 U217 ( .A1(n781), .A2(n576), .B1(n771), .B2(n578), .C1(n782), .C2(
        n86), .ZN(n769) );
  OAI222_X1 U218 ( .A1(n782), .A2(n90), .B1(n772), .B2(n91), .C1(n771), .C2(n4), .ZN(n770) );
  OAI222_X1 U219 ( .A1(n7560), .A2(n499), .B1(n743), .B2(n108), .C1(n7570), 
        .C2(n1), .ZN(n741) );
  OAI222_X1 U220 ( .A1(n7570), .A2(n107), .B1(n744), .B2(n501), .C1(n743), 
        .C2(n3), .ZN(n742) );
  NOR2_X1 U221 ( .A1(sub_64_I5_aco_B_0_), .A2(sub_64_I4_aco_B_0_), .ZN(n93) );
  NOR2_X1 U222 ( .A1(n67), .A2(sub_64_I8_aco_B_0_), .ZN(n464) );
  INV_X1 U223 ( .A(n695), .ZN(n344) );
  OAI222_X1 U224 ( .A1(n811), .A2(n423), .B1(n813), .B2(n424), .C1(n810), .C2(
        n425), .ZN(n695) );
  INV_X1 U225 ( .A(n696), .ZN(n343) );
  OAI222_X1 U226 ( .A1(n810), .A2(n423), .B1(n812), .B2(n424), .C1(n813), .C2(
        n425), .ZN(n696) );
  INV_X1 U227 ( .A(n646), .ZN(n298) );
  OAI222_X1 U228 ( .A1(n321), .A2(n401), .B1(n323), .B2(n402), .C1(n3200), 
        .C2(n403), .ZN(n646) );
  INV_X1 U229 ( .A(n647), .ZN(n297) );
  OAI222_X1 U230 ( .A1(n3200), .A2(n401), .B1(n322), .B2(n402), .C1(n323), 
        .C2(n403), .ZN(n647) );
  INV_X1 U231 ( .A(n672), .ZN(n321) );
  OAI222_X1 U232 ( .A1(n344), .A2(n411), .B1(n346), .B2(n412), .C1(n343), .C2(
        n413), .ZN(n672) );
  INV_X1 U233 ( .A(n673), .ZN(n3200) );
  OAI222_X1 U234 ( .A1(n343), .A2(n411), .B1(n345), .B2(n412), .C1(n346), .C2(
        n413), .ZN(n673) );
  CLKBUF_X1 U235 ( .A(n438), .Z(n122) );
  INV_X1 U236 ( .A(n718), .ZN(n811) );
  OAI222_X1 U237 ( .A1(n719), .A2(n122), .B1(n698), .B2(n440), .C1(n720), .C2(
        n442), .ZN(n718) );
  INV_X1 U238 ( .A(n7210), .ZN(n810) );
  OAI222_X1 U239 ( .A1(n720), .A2(n122), .B1(n699), .B2(n440), .C1(n698), .C2(
        n442), .ZN(n7210) );
  INV_X1 U240 ( .A(n5580), .ZN(n288) );
  OAI222_X1 U241 ( .A1(n312), .A2(n506), .B1(n3150), .B2(n4870), .C1(n3160), 
        .C2(n507), .ZN(n5580) );
  INV_X1 U242 ( .A(n560), .ZN(n3150) );
  INV_X1 U243 ( .A(n543), .ZN(n289) );
  OAI222_X1 U244 ( .A1(n3130), .A2(n506), .B1(n3160), .B2(n4870), .C1(n312), 
        .C2(n507), .ZN(n543) );
  INV_X1 U245 ( .A(n5210), .ZN(n290) );
  OAI222_X1 U246 ( .A1(n3140), .A2(n506), .B1(n312), .B2(n4870), .C1(n3130), 
        .C2(n507), .ZN(n5210) );
  INV_X1 U247 ( .A(n377), .ZN(n842) );
  INV_X1 U248 ( .A(n505), .ZN(n291) );
  OAI222_X1 U249 ( .A1(n311), .A2(n506), .B1(n3130), .B2(n4870), .C1(n3140), 
        .C2(n507), .ZN(n505) );
  INV_X1 U250 ( .A(n475), .ZN(n286) );
  OAI221_X1 U251 ( .B1(n299), .B2(n393), .C1(n287), .C2(n15), .A(n476), .ZN(
        n475) );
  INV_X1 U252 ( .A(n473), .ZN(n287) );
  AOI222_X1 U253 ( .A1(n125), .A2(n844), .B1(n846), .B2(n75), .C1(n845), .C2(
        n87), .ZN(n771) );
  AOI222_X1 U254 ( .A1(n7220), .A2(n121), .B1(n701), .B2(n466), .C1(n7230), 
        .C2(n468), .ZN(n698) );
  AOI222_X1 U255 ( .A1(n7580), .A2(n101), .B1(n745), .B2(n106), .C1(n7590), 
        .C2(n5), .ZN(n743) );
  OAI222_X1 U256 ( .A1(n771), .A2(n576), .B1(n7600), .B2(n578), .C1(n772), 
        .C2(n4), .ZN(n7580) );
  OAI222_X1 U257 ( .A1(n743), .A2(n499), .B1(n7240), .B2(n501), .C1(n744), 
        .C2(n3), .ZN(n7220) );
  INV_X1 U258 ( .A(n401), .ZN(n309) );
  INV_X1 U259 ( .A(n674), .ZN(n346) );
  OAI222_X1 U260 ( .A1(n813), .A2(n423), .B1(n815), .B2(n424), .C1(n812), .C2(
        n425), .ZN(n674) );
  INV_X1 U261 ( .A(n478), .ZN(n299) );
  OAI222_X1 U262 ( .A1(n325), .A2(n401), .B1(n334), .B2(n402), .C1(n324), .C2(
        n403), .ZN(n478) );
  INV_X1 U263 ( .A(n458), .ZN(n300) );
  OAI222_X1 U264 ( .A1(n326), .A2(n401), .B1(n324), .B2(n402), .C1(n325), .C2(
        n403), .ZN(n458) );
  INV_X1 U265 ( .A(n447), .ZN(n301) );
  OAI222_X1 U266 ( .A1(n327), .A2(n401), .B1(n325), .B2(n402), .C1(n326), .C2(
        n403), .ZN(n447) );
  INV_X1 U267 ( .A(n433), .ZN(n302) );
  OAI222_X1 U268 ( .A1(n328), .A2(n401), .B1(n326), .B2(n402), .C1(n327), .C2(
        n403), .ZN(n433) );
  INV_X1 U269 ( .A(n428), .ZN(n303) );
  OAI222_X1 U270 ( .A1(n329), .A2(n401), .B1(n327), .B2(n402), .C1(n328), .C2(
        n403), .ZN(n428) );
  INV_X1 U271 ( .A(n4200), .ZN(n304) );
  OAI222_X1 U272 ( .A1(n330), .A2(n401), .B1(n328), .B2(n402), .C1(n329), .C2(
        n403), .ZN(n4200) );
  INV_X1 U273 ( .A(n4160), .ZN(n305) );
  OAI222_X1 U274 ( .A1(n331), .A2(n401), .B1(n329), .B2(n402), .C1(n330), .C2(
        n403), .ZN(n4160) );
  INV_X1 U275 ( .A(n409), .ZN(n306) );
  OAI222_X1 U276 ( .A1(n332), .A2(n401), .B1(n330), .B2(n402), .C1(n331), .C2(
        n403), .ZN(n409) );
  INV_X1 U277 ( .A(n406), .ZN(n307) );
  OAI222_X1 U278 ( .A1(n322), .A2(n401), .B1(n331), .B2(n402), .C1(n332), .C2(
        n403), .ZN(n406) );
  INV_X1 U279 ( .A(n400), .ZN(n308) );
  OAI222_X1 U280 ( .A1(n323), .A2(n401), .B1(n332), .B2(n402), .C1(n322), .C2(
        n403), .ZN(n400) );
  INV_X1 U281 ( .A(n648), .ZN(n323) );
  OAI222_X1 U282 ( .A1(n346), .A2(n411), .B1(n3480), .B2(n412), .C1(n345), 
        .C2(n413), .ZN(n648) );
  CLKBUF_X1 U283 ( .A(n438), .Z(n123) );
  INV_X1 U284 ( .A(n697), .ZN(n813) );
  OAI222_X1 U285 ( .A1(n698), .A2(n123), .B1(n677), .B2(n440), .C1(n699), .C2(
        n442), .ZN(n697) );
  INV_X1 U286 ( .A(n613), .ZN(n292) );
  INV_X1 U287 ( .A(n5880), .ZN(n293) );
  INV_X1 U288 ( .A(n477), .ZN(n3101) );
  AOI222_X1 U289 ( .A1(n125), .A2(n845), .B1(n847), .B2(n75), .C1(n846), .C2(
        n87), .ZN(n772) );
  AOI222_X1 U290 ( .A1(n125), .A2(n846), .B1(n848), .B2(n75), .C1(n847), .C2(
        n89), .ZN(n7600) );
  AOI222_X1 U291 ( .A1(n7230), .A2(n120), .B1(n702), .B2(n466), .C1(n701), 
        .C2(n468), .ZN(n699) );
  AOI222_X1 U292 ( .A1(n701), .A2(n113), .B1(n680), .B2(n466), .C1(n702), .C2(
        n468), .ZN(n677) );
  AOI222_X1 U293 ( .A1(n7590), .A2(n100), .B1(n746), .B2(n104), .C1(n745), 
        .C2(n2), .ZN(n744) );
  AOI222_X1 U294 ( .A1(n745), .A2(n95), .B1(n7260), .B2(n105), .C1(n746), .C2(
        n2), .ZN(n7240) );
  OAI222_X1 U295 ( .A1(n772), .A2(n90), .B1(n7610), .B2(n91), .C1(n7600), .C2(
        n86), .ZN(n7590) );
  OAI222_X1 U296 ( .A1(n7600), .A2(n576), .B1(n747), .B2(n578), .C1(n7610), 
        .C2(n86), .ZN(n745) );
  OAI222_X1 U297 ( .A1(n744), .A2(n107), .B1(n7250), .B2(n109), .C1(n7240), 
        .C2(n1), .ZN(n7230) );
  OAI222_X1 U298 ( .A1(n7240), .A2(n499), .B1(n703), .B2(n109), .C1(n7250), 
        .C2(n1), .ZN(n701) );
  INV_X1 U299 ( .A(n493), .ZN(n324) );
  OAI222_X1 U300 ( .A1(n3500), .A2(n411), .B1(n806), .B2(n412), .C1(n3490), 
        .C2(n413), .ZN(n493) );
  INV_X1 U301 ( .A(n676), .ZN(n815) );
  OAI222_X1 U302 ( .A1(n677), .A2(n123), .B1(n6530), .B2(n440), .C1(n678), 
        .C2(n442), .ZN(n676) );
  INV_X1 U303 ( .A(n561), .ZN(n312) );
  OAI222_X1 U304 ( .A1(n337), .A2(n5230), .B1(n339), .B2(n508), .C1(n336), 
        .C2(n5240), .ZN(n561) );
  INV_X1 U305 ( .A(n563), .ZN(n339) );
  INV_X1 U306 ( .A(n544), .ZN(n3130) );
  OAI222_X1 U307 ( .A1(n338), .A2(n5230), .B1(n336), .B2(n508), .C1(n337), 
        .C2(n5240), .ZN(n544) );
  INV_X1 U308 ( .A(n675), .ZN(n345) );
  OAI222_X1 U309 ( .A1(n812), .A2(n423), .B1(n814), .B2(n424), .C1(n815), .C2(
        n425), .ZN(n675) );
  INV_X1 U310 ( .A(n650), .ZN(n3480) );
  OAI222_X1 U311 ( .A1(n815), .A2(n423), .B1(n817), .B2(n424), .C1(n814), .C2(
        n425), .ZN(n650) );
  INV_X1 U312 ( .A(n649), .ZN(n322) );
  OAI222_X1 U313 ( .A1(n345), .A2(n411), .B1(n3470), .B2(n412), .C1(n3480), 
        .C2(n413), .ZN(n649) );
  INV_X1 U314 ( .A(n479), .ZN(n325) );
  OAI222_X1 U315 ( .A1(n3510), .A2(n411), .B1(n3490), .B2(n412), .C1(n3500), 
        .C2(n413), .ZN(n479) );
  INV_X1 U316 ( .A(n459), .ZN(n326) );
  OAI222_X1 U317 ( .A1(n3520), .A2(n411), .B1(n3500), .B2(n412), .C1(n3510), 
        .C2(n413), .ZN(n459) );
  INV_X1 U318 ( .A(n448), .ZN(n327) );
  OAI222_X1 U319 ( .A1(n355), .A2(n411), .B1(n3510), .B2(n412), .C1(n3520), 
        .C2(n413), .ZN(n448) );
  INV_X1 U320 ( .A(n434), .ZN(n328) );
  OAI222_X1 U321 ( .A1(n503), .A2(n411), .B1(n3520), .B2(n412), .C1(n355), 
        .C2(n413), .ZN(n434) );
  INV_X1 U322 ( .A(n429), .ZN(n329) );
  OAI222_X1 U323 ( .A1(n541), .A2(n411), .B1(n355), .B2(n412), .C1(n503), .C2(
        n413), .ZN(n429) );
  INV_X1 U324 ( .A(n4210), .ZN(n330) );
  OAI222_X1 U325 ( .A1(n580), .A2(n411), .B1(n503), .B2(n412), .C1(n541), .C2(
        n413), .ZN(n4210) );
  INV_X1 U326 ( .A(n4170), .ZN(n331) );
  OAI222_X1 U327 ( .A1(n3470), .A2(n411), .B1(n541), .B2(n412), .C1(n580), 
        .C2(n413), .ZN(n4170) );
  INV_X1 U328 ( .A(n410), .ZN(n332) );
  OAI222_X1 U329 ( .A1(n3480), .A2(n411), .B1(n580), .B2(n412), .C1(n3470), 
        .C2(n413), .ZN(n410) );
  INV_X1 U330 ( .A(n700), .ZN(n812) );
  OAI222_X1 U331 ( .A1(n699), .A2(n122), .B1(n678), .B2(n440), .C1(n677), .C2(
        n442), .ZN(n700) );
  INV_X1 U332 ( .A(n5220), .ZN(n3140) );
  OAI222_X1 U333 ( .A1(n335), .A2(n5230), .B1(n337), .B2(n508), .C1(n338), 
        .C2(n5240), .ZN(n5220) );
  INV_X1 U334 ( .A(n5910), .ZN(n3160) );
  OAI221_X1 U335 ( .B1(n336), .B2(n5230), .C1(n5920), .C2(n78), .A(n593), .ZN(
        n5910) );
  INV_X1 U336 ( .A(n492), .ZN(n334) );
  INV_X1 U337 ( .A(n4890), .ZN(n311) );
  AOI222_X1 U338 ( .A1(n125), .A2(n847), .B1(n849), .B2(n69), .C1(n848), .C2(
        n88), .ZN(n7610) );
  AOI222_X1 U339 ( .A1(n702), .A2(n113), .B1(n681), .B2(n466), .C1(n680), .C2(
        n468), .ZN(n678) );
  AOI222_X1 U340 ( .A1(n746), .A2(n102), .B1(n7270), .B2(n106), .C1(n7260), 
        .C2(n5), .ZN(n7250) );
  OAI222_X1 U341 ( .A1(n7610), .A2(n90), .B1(n748), .B2(n91), .C1(n747), .C2(
        n4), .ZN(n746) );
  OAI222_X1 U342 ( .A1(n7250), .A2(n107), .B1(n704), .B2(n108), .C1(n703), 
        .C2(n3), .ZN(n702) );
  INV_X1 U343 ( .A(n679), .ZN(n814) );
  OAI222_X1 U344 ( .A1(n678), .A2(n123), .B1(n6540), .B2(n440), .C1(n6530), 
        .C2(n442), .ZN(n679) );
  INV_X1 U345 ( .A(n564), .ZN(n337) );
  OAI222_X1 U346 ( .A1(n525), .A2(n546), .B1(n565), .B2(n526), .C1(n547), .C2(
        n548), .ZN(n564) );
  INV_X1 U347 ( .A(n545), .ZN(n338) );
  OAI222_X1 U348 ( .A1(n528), .A2(n546), .B1(n547), .B2(n526), .C1(n525), .C2(
        n548), .ZN(n545) );
  INV_X1 U349 ( .A(n594), .ZN(n336) );
  OAI222_X1 U350 ( .A1(n547), .A2(n546), .B1(n526), .B2(n595), .C1(n565), .C2(
        n548), .ZN(n594) );
  OAI22_X1 U351 ( .A1(n548), .A2(n595), .B1(n565), .B2(n546), .ZN(n563) );
  NOR2_X1 U352 ( .A1(sub_64_I5_aco_B_0_), .A2(sub_64_I4_aco_B_0_), .ZN(n537)
         );
  INV_X1 U353 ( .A(n651), .ZN(n3470) );
  OAI222_X1 U354 ( .A1(n814), .A2(n423), .B1(n816), .B2(n424), .C1(n817), .C2(
        n425), .ZN(n651) );
  INV_X1 U355 ( .A(n514), .ZN(n3490) );
  OAI222_X1 U356 ( .A1(n819), .A2(n423), .B1(n8250), .B2(n424), .C1(n818), 
        .C2(n425), .ZN(n514) );
  INV_X1 U357 ( .A(n515), .ZN(n8250) );
  INV_X1 U358 ( .A(n513), .ZN(n806) );
  AOI222_X1 U359 ( .A1(n125), .A2(n848), .B1(n850), .B2(n70), .C1(n849), .C2(
        n87), .ZN(n747) );
  AOI222_X1 U360 ( .A1(n680), .A2(n115), .B1(n6560), .B2(n466), .C1(n681), 
        .C2(n468), .ZN(n6530) );
  AOI222_X1 U361 ( .A1(n681), .A2(n114), .B1(n6570), .B2(n466), .C1(n6560), 
        .C2(n468), .ZN(n6540) );
  AOI222_X1 U362 ( .A1(n7260), .A2(n102), .B1(n705), .B2(n104), .C1(n7270), 
        .C2(n5), .ZN(n703) );
  AOI222_X1 U363 ( .A1(n7270), .A2(n101), .B1(n706), .B2(n104), .C1(n705), 
        .C2(n2), .ZN(n704) );
  OAI222_X1 U364 ( .A1(n747), .A2(n576), .B1(n7280), .B2(n578), .C1(n748), 
        .C2(n4), .ZN(n7260) );
  OAI222_X1 U365 ( .A1(n748), .A2(n90), .B1(n729), .B2(n91), .C1(n7280), .C2(
        n86), .ZN(n7270) );
  OAI222_X1 U366 ( .A1(n703), .A2(n499), .B1(n682), .B2(n108), .C1(n704), .C2(
        n3), .ZN(n680) );
  OAI222_X1 U367 ( .A1(n704), .A2(n107), .B1(n683), .B2(n501), .C1(n682), .C2(
        n1), .ZN(n681) );
  AOI21_X1 U368 ( .B1(n76), .B2(n596), .A(n618), .ZN(n565) );
  NOR3_X1 U369 ( .A1(n76), .A2(n122), .A3(n6190), .ZN(n618) );
  AOI22_X1 U370 ( .A1(n76), .A2(n550), .B1(n566), .B2(sub_64_I12_aco_B_0_), 
        .ZN(n525) );
  AOI22_X1 U371 ( .A1(n596), .A2(sub_64_I12_aco_B_0_), .B1(n76), .B2(n566), 
        .ZN(n547) );
  AOI22_X1 U372 ( .A1(n76), .A2(n515), .B1(n550), .B2(sub_64_I12_aco_B_0_), 
        .ZN(n528) );
  INV_X1 U373 ( .A(n652), .ZN(n817) );
  OAI222_X1 U374 ( .A1(n6530), .A2(n124), .B1(n437), .B2(n440), .C1(n6540), 
        .C2(n442), .ZN(n652) );
  INV_X1 U375 ( .A(n6550), .ZN(n816) );
  OAI222_X1 U376 ( .A1(n6540), .A2(n124), .B1(n441), .B2(n440), .C1(n437), 
        .C2(n442), .ZN(n6550) );
  INV_X1 U377 ( .A(n494), .ZN(n3500) );
  OAI222_X1 U378 ( .A1(n820), .A2(n423), .B1(n818), .B2(n424), .C1(n819), .C2(
        n425), .ZN(n494) );
  INV_X1 U379 ( .A(n480), .ZN(n3510) );
  OAI222_X1 U380 ( .A1(n821), .A2(n423), .B1(n819), .B2(n424), .C1(n820), .C2(
        n425), .ZN(n480) );
  INV_X1 U381 ( .A(n460), .ZN(n3520) );
  OAI222_X1 U382 ( .A1(n822), .A2(n423), .B1(n820), .B2(n424), .C1(n821), .C2(
        n425), .ZN(n460) );
  INV_X1 U383 ( .A(n4490), .ZN(n355) );
  OAI222_X1 U384 ( .A1(n8230), .A2(n423), .B1(n821), .B2(n424), .C1(n822), 
        .C2(n425), .ZN(n4490) );
  INV_X1 U385 ( .A(n435), .ZN(n503) );
  OAI222_X1 U386 ( .A1(n8240), .A2(n423), .B1(n822), .B2(n424), .C1(n8230), 
        .C2(n425), .ZN(n435) );
  INV_X1 U387 ( .A(n430), .ZN(n541) );
  OAI222_X1 U388 ( .A1(n816), .A2(n423), .B1(n8230), .B2(n424), .C1(n8240), 
        .C2(n425), .ZN(n430) );
  INV_X1 U389 ( .A(n4220), .ZN(n580) );
  OAI222_X1 U390 ( .A1(n817), .A2(n423), .B1(n8240), .B2(n424), .C1(n816), 
        .C2(n425), .ZN(n4220) );
  AOI222_X1 U391 ( .A1(n6560), .A2(n119), .B1(n463), .B2(n466), .C1(n6570), 
        .C2(n468), .ZN(n437) );
  AOI222_X1 U392 ( .A1(n705), .A2(n98), .B1(n684), .B2(n105), .C1(n706), .C2(
        n2), .ZN(n682) );
  OAI222_X1 U393 ( .A1(n7280), .A2(n576), .B1(n707), .B2(n578), .C1(n729), 
        .C2(n86), .ZN(n705) );
  OAI222_X1 U394 ( .A1(n682), .A2(n499), .B1(n6580), .B2(n501), .C1(n683), 
        .C2(n1), .ZN(n6560) );
  INV_X1 U395 ( .A(n532), .ZN(n818) );
  OAI222_X1 U396 ( .A1(n496), .A2(n124), .B1(n533), .B2(n440), .C1(n5170), 
        .C2(n442), .ZN(n532) );
  INV_X1 U397 ( .A(n516), .ZN(n819) );
  OAI222_X1 U398 ( .A1(n482), .A2(n122), .B1(n5170), .B2(n440), .C1(n496), 
        .C2(n442), .ZN(n516) );
  INV_X1 U399 ( .A(n495), .ZN(n820) );
  OAI222_X1 U400 ( .A1(n462), .A2(n122), .B1(n496), .B2(n440), .C1(n482), .C2(
        n442), .ZN(n495) );
  INV_X1 U401 ( .A(n481), .ZN(n821) );
  OAI222_X1 U402 ( .A1(n4510), .A2(n122), .B1(n482), .B2(n440), .C1(n462), 
        .C2(n442), .ZN(n481) );
  INV_X1 U403 ( .A(n461), .ZN(n822) );
  OAI222_X1 U404 ( .A1(n439), .A2(n123), .B1(n462), .B2(n440), .C1(n4510), 
        .C2(n442), .ZN(n461) );
  INV_X1 U405 ( .A(n4500), .ZN(n8230) );
  OAI222_X1 U406 ( .A1(n441), .A2(n123), .B1(n4510), .B2(n440), .C1(n439), 
        .C2(n442), .ZN(n4500) );
  INV_X1 U407 ( .A(n436), .ZN(n8240) );
  OAI222_X1 U408 ( .A1(n437), .A2(n123), .B1(n439), .B2(n440), .C1(n441), .C2(
        n442), .ZN(n436) );
  OAI22_X1 U409 ( .A1(sub_64_I11_aco_B_0_), .A2(n5510), .B1(n567), .B2(n5520), 
        .ZN(n550) );
  OAI21_X1 U410 ( .B1(sub_64_I11_aco_B_0_), .B2(n597), .A(n6200), .ZN(n596) );
  NAND3_X1 U411 ( .A1(sub_64_I11_aco_B_0_), .A2(n83), .A3(n8270), .ZN(n6200)
         );
  INV_X1 U412 ( .A(n3830), .ZN(n849) );
  OR3_X1 U413 ( .A1(n123), .A2(sub_64_I12_aco_B_0_), .A3(n6190), .ZN(n595) );
  AOI222_X1 U414 ( .A1(n497), .A2(n113), .B1(n534), .B2(n466), .C1(n5180), 
        .C2(n468), .ZN(n496) );
  AOI222_X1 U415 ( .A1(n4830), .A2(n113), .B1(n5180), .B2(n466), .C1(n497), 
        .C2(n468), .ZN(n482) );
  AOI222_X1 U416 ( .A1(n6570), .A2(n118), .B1(n467), .B2(n466), .C1(n463), 
        .C2(n468), .ZN(n441) );
  AOI222_X1 U417 ( .A1(n465), .A2(n113), .B1(n497), .B2(n466), .C1(n4830), 
        .C2(n468), .ZN(n462) );
  AOI222_X1 U418 ( .A1(n467), .A2(n113), .B1(n4830), .B2(n466), .C1(n465), 
        .C2(n468), .ZN(n4510) );
  AOI222_X1 U419 ( .A1(n463), .A2(n113), .B1(n465), .B2(n466), .C1(n467), .C2(
        n468), .ZN(n439) );
  AOI222_X1 U420 ( .A1(n706), .A2(n100), .B1(n685), .B2(n106), .C1(n684), .C2(
        n5), .ZN(n683) );
  AOI222_X1 U421 ( .A1(n5180), .A2(n113), .B1(n5540), .B2(n466), .C1(n534), 
        .C2(n468), .ZN(n5170) );
  OAI222_X1 U422 ( .A1(n729), .A2(n90), .B1(n708), .B2(n91), .C1(n707), .C2(n4), .ZN(n706) );
  OAI222_X1 U423 ( .A1(n683), .A2(n107), .B1(n6590), .B2(n109), .C1(n6580), 
        .C2(n3), .ZN(n6570) );
  OAI222_X1 U424 ( .A1(n6580), .A2(n499), .B1(n498), .B2(n109), .C1(n6590), 
        .C2(n3), .ZN(n463) );
  OAI21_X1 U425 ( .B1(n67), .B2(n599), .A(n6210), .ZN(n598) );
  NAND3_X1 U426 ( .A1(n67), .A2(n77), .A3(n6220), .ZN(n6210) );
  INV_X1 U427 ( .A(n3810), .ZN(n850) );
  INV_X1 U428 ( .A(n3820), .ZN(n851) );
  INV_X1 U429 ( .A(n533), .ZN(n8260) );
  AOI222_X1 U430 ( .A1(n125), .A2(n853), .B1(n855), .B2(n75), .C1(n854), .C2(
        n89), .ZN(n708) );
  AOI222_X1 U431 ( .A1(n684), .A2(n103), .B1(n6600), .B2(n104), .C1(n685), 
        .C2(n5), .ZN(n6580) );
  AOI222_X1 U432 ( .A1(n685), .A2(n103), .B1(n661), .B2(n105), .C1(n6600), 
        .C2(n2), .ZN(n6590) );
  OAI222_X1 U433 ( .A1(n707), .A2(n576), .B1(n686), .B2(n578), .C1(n708), .C2(
        n4), .ZN(n684) );
  OAI222_X1 U434 ( .A1(n708), .A2(n90), .B1(n6870), .B2(n91), .C1(n686), .C2(
        n86), .ZN(n685) );
  OAI222_X1 U435 ( .A1(n535), .A2(n107), .B1(n831), .B2(n501), .C1(n5550), 
        .C2(n3), .ZN(n534) );
  INV_X1 U436 ( .A(n573), .ZN(n831) );
  OAI222_X1 U437 ( .A1(n6590), .A2(n107), .B1(n502), .B2(n108), .C1(n498), 
        .C2(n1), .ZN(n467) );
  INV_X1 U438 ( .A(n374), .ZN(n852) );
  AOI222_X1 U439 ( .A1(n125), .A2(n854), .B1(n856), .B2(n75), .C1(n855), .C2(
        n88), .ZN(n686) );
  AOI222_X1 U440 ( .A1(n125), .A2(n855), .B1(n8570), .B2(n75), .C1(n856), .C2(
        n87), .ZN(n6870) );
  AOI222_X1 U441 ( .A1(n6600), .A2(n94), .B1(n536), .B2(n106), .C1(n661), .C2(
        n2), .ZN(n498) );
  OAI222_X1 U442 ( .A1(n686), .A2(n576), .B1(n662), .B2(n578), .C1(n6870), 
        .C2(n86), .ZN(n6600) );
  OAI222_X1 U443 ( .A1(n5190), .A2(n499), .B1(n5550), .B2(n108), .C1(n535), 
        .C2(n1), .ZN(n5180) );
  OAI222_X1 U444 ( .A1(n500), .A2(n107), .B1(n535), .B2(n109), .C1(n5190), 
        .C2(n1), .ZN(n497) );
  OAI222_X1 U445 ( .A1(n502), .A2(n107), .B1(n5190), .B2(n501), .C1(n500), 
        .C2(n3), .ZN(n4830) );
  OAI222_X1 U446 ( .A1(n498), .A2(n499), .B1(n500), .B2(n108), .C1(n502), .C2(
        n3), .ZN(n465) );
  INV_X1 U447 ( .A(n372), .ZN(n853) );
  AOI222_X1 U448 ( .A1(n125), .A2(n856), .B1(n8580), .B2(n69), .C1(n8570), 
        .C2(n88), .ZN(n662) );
  AOI222_X1 U449 ( .A1(n538), .A2(n95), .B1(n574), .B2(n105), .C1(n5560), .C2(
        n2), .ZN(n535) );
  AOI222_X1 U450 ( .A1(n540), .A2(n96), .B1(n5560), .B2(n104), .C1(n538), .C2(
        n5), .ZN(n5190) );
  AOI222_X1 U451 ( .A1(n536), .A2(n970), .B1(n538), .B2(n104), .C1(n540), .C2(
        n5), .ZN(n500) );
  AOI222_X1 U452 ( .A1(n661), .A2(n94), .B1(n540), .B2(n106), .C1(n536), .C2(
        n5), .ZN(n502) );
  OAI222_X1 U453 ( .A1(n6870), .A2(n90), .B1(n663), .B2(n91), .C1(n662), .C2(
        n4), .ZN(n661) );
  OAI222_X1 U454 ( .A1(n662), .A2(n90), .B1(n575), .B2(n578), .C1(n663), .C2(
        n4), .ZN(n536) );
  OAI21_X1 U455 ( .B1(sub_64_I5_aco_B_0_), .B2(n607), .A(n627), .ZN(n573) );
  NAND3_X1 U456 ( .A1(sub_64_I5_aco_B_0_), .A2(n628), .A3(n6260), .ZN(n627) );
  AOI22_X1 U457 ( .A1(n628), .A2(n574), .B1(sub_64_I4_aco_B_0_), .B2(n6260), 
        .ZN(n607) );
  INV_X1 U458 ( .A(n373), .ZN(n854) );
  AOI222_X1 U459 ( .A1(n125), .A2(n8570), .B1(n8590), .B2(n70), .C1(n8580), 
        .C2(n89), .ZN(n663) );
  OAI222_X1 U460 ( .A1(n663), .A2(n90), .B1(n579), .B2(n91), .C1(n575), .C2(
        n86), .ZN(n540) );
  OAI222_X1 U461 ( .A1(n575), .A2(n576), .B1(n577), .B2(n91), .C1(n579), .C2(
        n4), .ZN(n538) );
  NOR2_X1 U462 ( .A1(n631), .A2(n90), .ZN(n6260) );
  AOI222_X1 U463 ( .A1(n125), .A2(n8590), .B1(n8610), .B2(n73), .C1(n8600), 
        .C2(n87), .ZN(n579) );
  INV_X1 U464 ( .A(n371), .ZN(n8610) );
  AOI221_X1 U465 ( .B1(n125), .B2(n8600), .C1(n632), .C2(n75), .A(n633), .ZN(
        n577) );
  NOR3_X1 U466 ( .A1(n74), .A2(n125), .A3(n371), .ZN(n633) );
  INV_X1 U467 ( .A(n369), .ZN(n8580) );
  INV_X1 U468 ( .A(n367), .ZN(n8590) );
  INV_X1 U469 ( .A(n368), .ZN(n8600) );
  NAND4_X1 U470 ( .A1(n376), .A2(n377), .A3(n378), .A4(n379), .ZN(n363) );
  NOR4_X1 U471 ( .A1(n380), .A2(n846), .A3(n848), .A4(n847), .ZN(n379) );
  NOR3_X1 U472 ( .A1(n843), .A2(n845), .A3(n844), .ZN(n378) );
  NAND3_X1 U473 ( .A1(n3810), .A2(n3820), .A3(n3830), .ZN(n380) );
  NOR3_X1 U474 ( .A1(n855), .A2(n8570), .A3(n856), .ZN(n375) );
  NOR4_X1 U475 ( .A1(N226), .A2(N225), .A3(N224), .A4(n128), .ZN(n803) );
  XNOR2_X1 U476 ( .A(n147), .B(a[23]), .ZN(shamt[0]) );
  BUF_X1 U477 ( .A(n141), .Z(n146) );
  INV_X1 U478 ( .A(a[23]), .ZN(n14) );
  NOR3_X1 U479 ( .A1(N229), .A2(N231), .A3(N230), .ZN(n802) );
  OR2_X1 U480 ( .A1(add_42_B_0_), .A2(a[23]), .ZN(sub_46_ni_carry[1]) );
  OR2_X1 U481 ( .A1(n603), .A2(N483), .ZN(sub_64_I7_aco_carry[1]) );
  OR2_X1 U482 ( .A1(n606), .A2(N415), .ZN(sub_64_I5_aco_carry[1]) );
  OR2_X1 U483 ( .A1(n571), .A2(N551), .ZN(sub_64_I9_aco_carry[1]) );
  OR2_X1 U484 ( .A1(n5520), .A2(N619), .ZN(sub_64_I11_aco_carry[1]) );
  OR2_X1 U485 ( .A1(n530), .A2(N687), .ZN(sub_64_I13_aco_carry[1]) );
  OR2_X1 U486 ( .A1(n4900), .A2(N823), .ZN(sub_64_I17_aco_carry[1]) );
  OR2_X1 U487 ( .A1(n511), .A2(N755), .ZN(sub_64_I15_aco_carry[1]) );
  OR2_X1 U488 ( .A1(a[27]), .A2(sub_46_ni_carry[4]), .ZN(sub_46_ni_carry[5])
         );
  OR2_X1 U489 ( .A1(a[26]), .A2(sub_46_ni_carry[3]), .ZN(sub_46_ni_carry[4])
         );
  OR2_X1 U490 ( .A1(a[25]), .A2(sub_46_ni_carry[2]), .ZN(sub_46_ni_carry[3])
         );
  OR2_X1 U491 ( .A1(a[24]), .A2(sub_46_ni_carry[1]), .ZN(sub_46_ni_carry[2])
         );
  NAND2_X1 U492 ( .A1(n511), .A2(n82), .ZN(n411) );
  INV_X1 U493 ( .A(n139), .ZN(n129) );
  XNOR2_X1 U494 ( .A(n474), .B(N891), .ZN(N925) );
  XNOR2_X1 U495 ( .A(n630), .B(N313), .ZN(N347) );
  XNOR2_X1 U496 ( .A(n568), .B(N585), .ZN(N619) );
  XNOR2_X1 U497 ( .A(n6240), .B(N449), .ZN(N483) );
  XNOR2_X1 U498 ( .A(n562), .B(N789), .ZN(N823) );
  XNOR2_X1 U499 ( .A(n549), .B(N653), .ZN(N687) );
  XNOR2_X1 U500 ( .A(n529), .B(N721), .ZN(N755) );
  XNOR2_X1 U501 ( .A(n457), .B(N925), .ZN(N959) );
  XNOR2_X1 U502 ( .A(n628), .B(N381), .ZN(N415) );
  XNOR2_X1 U503 ( .A(n600), .B(N517), .ZN(N551) );
  XNOR2_X1 U504 ( .A(n5520), .B(N619), .ZN(N653) );
  XNOR2_X1 U505 ( .A(n603), .B(N483), .ZN(N517) );
  XNOR2_X1 U506 ( .A(n4900), .B(N823), .ZN(N857) );
  XNOR2_X1 U507 ( .A(n511), .B(N755), .ZN(N789) );
  XNOR2_X1 U508 ( .A(n530), .B(N687), .ZN(N721) );
  XNOR2_X1 U509 ( .A(n606), .B(N415), .ZN(N449) );
  XNOR2_X1 U510 ( .A(n571), .B(N551), .ZN(N585) );
  XNOR2_X1 U511 ( .A(n125), .B(a[23]), .ZN(N224) );
  AOI22_X1 U512 ( .A1(N186), .A2(n129), .B1(N221), .B2(n137), .ZN(n376) );
  XNOR2_X1 U513 ( .A(a[24]), .B(sub_46_ni_carry[1]), .ZN(N225) );
  XNOR2_X1 U514 ( .A(a[25]), .B(sub_46_ni_carry[2]), .ZN(N226) );
  XNOR2_X1 U515 ( .A(sub_64_aco_A_1_), .B(sub_64_aco_carry[1]), .ZN(N314) );
  OAI221_X1 U516 ( .B1(n270), .B2(n4520), .C1(n443), .C2(n3840), .A(n4530), 
        .ZN(out[9]) );
  XOR2_X1 U517 ( .A(a[26]), .B(sub_46_ni_carry[3]), .Z(n8) );
  INV_X1 U518 ( .A(n360), .ZN(sub_64_aco_A_0_) );
  AOI22_X1 U519 ( .A1(n138), .A2(N224), .B1(n128), .B2(n7), .ZN(n360) );
  INV_X1 U520 ( .A(n370), .ZN(n840) );
  XOR2_X1 U521 ( .A(a[27]), .B(sub_46_ni_carry[4]), .Z(n9) );
  AND2_X1 U522 ( .A1(Out_Exponent[0]), .A2(n837), .ZN(out[23]) );
  XNOR2_X1 U523 ( .A(n582), .B(N993), .ZN(Out_Exponent[0]) );
  INV_X1 U524 ( .A(n138), .ZN(n128) );
  AOI22_X1 U525 ( .A1(N185), .A2(n129), .B1(N220), .B2(n136), .ZN(n377) );
  INV_X1 U526 ( .A(n804), .ZN(n843) );
  AOI22_X1 U527 ( .A1(N184), .A2(n129), .B1(N219), .B2(n137), .ZN(n804) );
  OAI221_X1 U528 ( .B1(n3140), .B2(n4870), .C1(n63), .C2(n3101), .A(n4880), 
        .ZN(n473) );
  INV_X1 U529 ( .A(n7920), .ZN(n844) );
  AOI22_X1 U530 ( .A1(N183), .A2(n129), .B1(N218), .B2(n136), .ZN(n7920) );
  INV_X1 U531 ( .A(n7930), .ZN(n845) );
  AOI22_X1 U532 ( .A1(N182), .A2(n129), .B1(N217), .B2(n134), .ZN(n7930) );
  OAI221_X1 U533 ( .B1(n338), .B2(n508), .C1(sub_64_I16_aco_B_0_), .C2(n334), 
        .A(n509), .ZN(n4890) );
  INV_X1 U534 ( .A(n784), .ZN(n847) );
  AOI22_X1 U535 ( .A1(N180), .A2(n129), .B1(N215), .B2(n135), .ZN(n784) );
  INV_X1 U536 ( .A(n783), .ZN(n846) );
  AOI22_X1 U537 ( .A1(N181), .A2(n129), .B1(N216), .B2(n135), .ZN(n783) );
  INV_X1 U538 ( .A(n773), .ZN(n848) );
  AOI22_X1 U539 ( .A1(N179), .A2(n129), .B1(N214), .B2(n134), .ZN(n773) );
  AOI22_X1 U540 ( .A1(N178), .A2(n129), .B1(N213), .B2(n135), .ZN(n3830) );
  AOI221_X1 U541 ( .B1(n534), .B2(n113), .C1(n8280), .C2(n67), .A(n570), .ZN(
        n533) );
  INV_X1 U542 ( .A(n572), .ZN(n8280) );
  AOI22_X1 U543 ( .A1(N176), .A2(n129), .B1(N211), .B2(n134), .ZN(n3820) );
  AOI22_X1 U544 ( .A1(N177), .A2(n128), .B1(N212), .B2(n133), .ZN(n3810) );
  AOI22_X1 U545 ( .A1(N175), .A2(n128), .B1(N210), .B2(n133), .ZN(n374) );
  AOI22_X1 U546 ( .A1(N174), .A2(n128), .B1(N209), .B2(n133), .ZN(n372) );
  AND3_X1 U547 ( .A1(sub_64_I6_aco_B_0_), .A2(n103), .A3(n6260), .ZN(n6250) );
  AOI221_X1 U548 ( .B1(n5560), .B2(n94), .C1(n832), .C2(sub_64_I5_aco_B_0_), 
        .A(n605), .ZN(n5550) );
  INV_X1 U549 ( .A(n607), .ZN(n832) );
  AOI22_X1 U550 ( .A1(N173), .A2(n128), .B1(N208), .B2(n132), .ZN(n373) );
  INV_X1 U551 ( .A(n730), .ZN(n855) );
  AOI22_X1 U552 ( .A1(N172), .A2(n128), .B1(N207), .B2(n132), .ZN(n730) );
  INV_X1 U553 ( .A(n709), .ZN(n856) );
  AOI22_X1 U554 ( .A1(N171), .A2(n128), .B1(N206), .B2(n132), .ZN(n709) );
  INV_X1 U555 ( .A(n710), .ZN(n8570) );
  AOI22_X1 U556 ( .A1(N170), .A2(n128), .B1(N205), .B2(n131), .ZN(n710) );
  AOI22_X1 U557 ( .A1(N169), .A2(n128), .B1(N204), .B2(n131), .ZN(n369) );
  AOI22_X1 U558 ( .A1(N168), .A2(n128), .B1(N203), .B2(n131), .ZN(n367) );
  AOI22_X1 U559 ( .A1(N167), .A2(n128), .B1(N202), .B2(n130), .ZN(n368) );
  AOI22_X1 U560 ( .A1(N166), .A2(n128), .B1(N201), .B2(n130), .ZN(n371) );
  OAI211_X1 U561 ( .C1(n140), .C2(n8620), .A(n370), .B(n371), .ZN(n365) );
  INV_X1 U562 ( .A(N165), .ZN(n8620) );
  OR4_X1 U563 ( .A1(N586), .A2(N585), .A3(N588), .A4(N587), .ZN(n752) );
  OR4_X1 U564 ( .A1(N654), .A2(N653), .A3(N656), .A4(N655), .ZN(n734) );
  OR4_X1 U565 ( .A1(N790), .A2(N789), .A3(N792), .A4(N791), .ZN(n6910) );
  OR4_X1 U566 ( .A1(N722), .A2(N721), .A3(N724), .A4(N723), .ZN(n714) );
  OR4_X1 U567 ( .A1(N926), .A2(N925), .A3(N928), .A4(N927), .ZN(n642) );
  OR4_X1 U568 ( .A1(N314), .A2(N313), .A3(N316), .A4(N315), .ZN(n797) );
  OR4_X1 U570 ( .A1(N382), .A2(N381), .A3(N384), .A4(N383), .ZN(n788) );
  OR4_X1 U571 ( .A1(N518), .A2(N517), .A3(N520), .A4(N519), .ZN(n765) );
  OAI22_X1 U572 ( .A1(n32), .A2(n228), .B1(n60), .B2(n871), .ZN(inShift[7]) );
  OAI22_X1 U573 ( .A1(n24), .A2(n8920), .B1(n144), .B2(n238), .ZN(inShift[6])
         );
  OAI22_X1 U574 ( .A1(n53), .A2(n8930), .B1(n145), .B2(n237), .ZN(inShift[4])
         );
  OAI22_X1 U575 ( .A1(n3100), .A2(n227), .B1(n54), .B2(n872), .ZN(inShift[5])
         );
  OAI22_X1 U576 ( .A1(n37), .A2(n8910), .B1(n54), .B2(n239), .ZN(inShift[8])
         );
  OAI22_X1 U577 ( .A1(n34), .A2(n2260), .B1(n65), .B2(n873), .ZN(inShift[3])
         );
  OAI22_X1 U578 ( .A1(n45), .A2(n2250), .B1(n60), .B2(n874), .ZN(inShift[2])
         );
  OAI22_X1 U579 ( .A1(n27), .A2(n886), .B1(n64), .B2(n244), .ZN(inShift[18])
         );
  OAI22_X1 U580 ( .A1(n25), .A2(n2310), .B1(n65), .B2(n868), .ZN(inShift[13])
         );
  OAI22_X1 U581 ( .A1(n28), .A2(n890), .B1(n59), .B2(n240), .ZN(inShift[10])
         );
  OAI22_X1 U582 ( .A1(n52), .A2(n889), .B1(n57), .B2(n241), .ZN(inShift[12])
         );
  OAI22_X1 U583 ( .A1(n33), .A2(n885), .B1(n60), .B2(n865), .ZN(inShift[19])
         );
  OAI22_X1 U584 ( .A1(n43), .A2(n234), .B1(n60), .B2(n8640), .ZN(inShift[21])
         );
  OAI22_X1 U585 ( .A1(n49), .A2(n2300), .B1(n55), .B2(n869), .ZN(inShift[11])
         );
  XNOR2_X1 U586 ( .A(a[29]), .B(sub_46_ni_carry[6]), .ZN(N230) );
  XNOR2_X1 U587 ( .A(a[28]), .B(sub_46_ni_carry[5]), .ZN(N229) );
  OAI22_X1 U588 ( .A1(n23), .A2(n884), .B1(n61), .B2(n245), .ZN(inShift[20])
         );
  OAI22_X1 U589 ( .A1(n30), .A2(n887), .B1(n61), .B2(n243), .ZN(inShift[16])
         );
  OAI22_X1 U590 ( .A1(n47), .A2(n888), .B1(n61), .B2(n242), .ZN(inShift[14])
         );
  OAI22_X1 U591 ( .A1(n51), .A2(n232), .B1(n59), .B2(n867), .ZN(inShift[15])
         );
  XNOR2_X1 U592 ( .A(N966), .B(sub_64_I21_aco_carry[7]), .ZN(N1000) );
  XNOR2_X1 U593 ( .A(N558), .B(sub_64_I9_aco_carry[7]), .ZN(N592) );
  XNOR2_X1 U594 ( .A(N626), .B(sub_64_I11_aco_carry[7]), .ZN(N660) );
  XNOR2_X1 U595 ( .A(N694), .B(sub_64_I13_aco_carry[7]), .ZN(N728) );
  XNOR2_X1 U596 ( .A(N898), .B(sub_64_I19_aco_carry[7]), .ZN(N932) );
  XNOR2_X1 U597 ( .A(N762), .B(sub_64_I15_aco_carry[7]), .ZN(N796) );
  XNOR2_X1 U598 ( .A(N864), .B(sub_64_I18_aco_carry[7]), .ZN(N898) );
  XNOR2_X1 U599 ( .A(N932), .B(sub_64_I20_aco_carry[7]), .ZN(N966) );
  XOR2_X1 U600 ( .A(n3540), .B(sub_64_aco_carry[7]), .Z(N320) );
  AOI22_X1 U601 ( .A1(n137), .A2(N231), .B1(n128), .B2(N198), .ZN(n3540) );
  XNOR2_X1 U602 ( .A(N354), .B(sub_64_I3_aco_carry[7]), .ZN(N388) );
  XNOR2_X1 U603 ( .A(N524), .B(sub_64_I8_aco_carry[7]), .ZN(N558) );
  XNOR2_X1 U604 ( .A(N422), .B(sub_64_I5_aco_carry[7]), .ZN(N456) );
  XNOR2_X1 U605 ( .A(N320), .B(sub_64_I2_aco_carry[7]), .ZN(N354) );
  XNOR2_X1 U606 ( .A(N592), .B(sub_64_I10_aco_carry[7]), .ZN(N626) );
  XNOR2_X1 U607 ( .A(N490), .B(sub_64_I7_aco_carry[7]), .ZN(N524) );
  XNOR2_X1 U608 ( .A(N388), .B(sub_64_I4_aco_carry[7]), .ZN(N422) );
  XNOR2_X1 U609 ( .A(N660), .B(sub_64_I12_aco_carry[7]), .ZN(N694) );
  XNOR2_X1 U610 ( .A(N456), .B(sub_64_I6_aco_carry[7]), .ZN(N490) );
  XNOR2_X1 U611 ( .A(N728), .B(sub_64_I14_aco_carry[7]), .ZN(N762) );
  XNOR2_X1 U612 ( .A(N830), .B(sub_64_I17_aco_carry[7]), .ZN(N864) );
  XNOR2_X1 U613 ( .A(N796), .B(sub_64_I16_aco_carry[7]), .ZN(N830) );
  OR4_X1 U614 ( .A1(N450), .A2(N449), .A3(N452), .A4(N451), .ZN(n777) );
  INV_X1 U615 ( .A(b[25]), .ZN(n149) );
  NAND2_X1 U616 ( .A1(b[23]), .A2(n14), .ZN(sub_36_carry[1]) );
  BUF_X1 U617 ( .A(n3530), .Z(n21) );
  INV_X1 U618 ( .A(b[26]), .ZN(n150) );
  INV_X1 U619 ( .A(n754), .ZN(n8290) );
  INV_X1 U620 ( .A(b[27]), .ZN(n151) );
  OAI22_X1 U621 ( .A1(n36), .A2(n878), .B1(n145), .B2(n1980), .ZN(b[27]) );
  OAI221_X2 U622 ( .B1(n785), .B2(n786), .C1(n833), .C2(n628), .A(n834), .ZN(
        n606) );
  INV_X1 U623 ( .A(n779), .ZN(n833) );
  BUF_X1 U624 ( .A(n20), .Z(n141) );
  OAI22_X1 U625 ( .A1(n48), .A2(n2240), .B1(n60), .B2(n875), .ZN(inShift[1])
         );
  OAI221_X2 U626 ( .B1(n639), .B2(n640), .C1(n273), .C2(n80), .A(n274), .ZN(
        n4550) );
  XNOR2_X1 U627 ( .A(a[30]), .B(sub_46_ni_carry[7]), .ZN(N231) );
  NAND2_X1 U628 ( .A1(n12), .A2(n13), .ZN(sub_46_ni_carry[7]) );
  INV_X1 U629 ( .A(a[29]), .ZN(n12) );
  INV_X1 U630 ( .A(sub_46_ni_carry[6]), .ZN(n13) );
  OAI22_X1 U631 ( .A1(n35), .A2(n8940), .B1(n144), .B2(n235), .ZN(inShift[0])
         );
  XNOR2_X1 U632 ( .A(N1000), .B(sub_64_I22_aco_carry[7]), .ZN(Out_Exponent[7])
         );
  AND2_X1 U633 ( .A1(Out_Exponent[5]), .A2(n837), .ZN(out[28]) );
  AND2_X1 U634 ( .A1(Out_Exponent[4]), .A2(n837), .ZN(out[27]) );
  OAI22_X1 U635 ( .A1(n146), .A2(n241), .B1(n64), .B2(n889), .ZN(a[12]) );
  OAI22_X1 U636 ( .A1(n25), .A2(n242), .B1(n65), .B2(n888), .ZN(a[14]) );
  OAI22_X1 U637 ( .A1(n21), .A2(n240), .B1(n60), .B2(n890), .ZN(a[10]) );
  OAI22_X1 U638 ( .A1(n141), .A2(n869), .B1(n61), .B2(n2300), .ZN(a[11]) );
  OAI22_X1 U639 ( .A1(n53), .A2(n244), .B1(n61), .B2(n886), .ZN(a[18]) );
  OAI22_X1 U640 ( .A1(n24), .A2(n243), .B1(n145), .B2(n887), .ZN(a[16]) );
  OAI22_X1 U641 ( .A1(n34), .A2(n866), .B1(n144), .B2(n233), .ZN(a[17]) );
  OAI22_X1 U642 ( .A1(n26), .A2(n868), .B1(n59), .B2(n2310), .ZN(a[13]) );
  OAI22_X1 U643 ( .A1(n23), .A2(n867), .B1(n143), .B2(n232), .ZN(a[15]) );
  NOR4_X1 U644 ( .A1(N193), .A2(N192), .A3(n7), .A4(n130), .ZN(n801) );
  XNOR2_X1 U645 ( .A(N348), .B(sub_64_I3_aco_carry[1]), .ZN(N382) );
  XNOR2_X1 U646 ( .A(N416), .B(sub_64_I5_aco_carry[1]), .ZN(N450) );
  XNOR2_X1 U647 ( .A(N484), .B(sub_64_I7_aco_carry[1]), .ZN(N518) );
  XNOR2_X1 U648 ( .A(N824), .B(sub_64_I17_aco_carry[1]), .ZN(N858) );
  XNOR2_X1 U649 ( .A(N552), .B(sub_64_I9_aco_carry[1]), .ZN(N586) );
  XNOR2_X1 U650 ( .A(N620), .B(sub_64_I11_aco_carry[1]), .ZN(N654) );
  XNOR2_X1 U651 ( .A(N756), .B(sub_64_I15_aco_carry[1]), .ZN(N790) );
  XNOR2_X1 U652 ( .A(N688), .B(sub_64_I13_aco_carry[1]), .ZN(N722) );
  XNOR2_X1 U653 ( .A(N960), .B(sub_64_I21_aco_carry[1]), .ZN(N994) );
  BUF_X1 U654 ( .A(n6), .Z(n139) );
  OAI22_X1 U655 ( .A1(n41), .A2(n235), .B1(n60), .B2(n8940), .ZN(a[0]) );
  OAI22_X1 U656 ( .A1(n42), .A2(n883), .B1(n64), .B2(n246), .ZN(inShift[22])
         );
  INV_X1 U657 ( .A(n359), .ZN(sub_64_aco_A_1_) );
  AOI22_X1 U658 ( .A1(n138), .A2(N225), .B1(n128), .B2(N192), .ZN(n359) );
  INV_X1 U659 ( .A(N195), .ZN(n838) );
  INV_X1 U660 ( .A(N194), .ZN(n839) );
  AND2_X1 U661 ( .A1(Out_Exponent[3]), .A2(n837), .ZN(out[26]) );
  AND2_X1 U662 ( .A1(Out_Exponent[2]), .A2(n837), .ZN(out[25]) );
  AND2_X1 U663 ( .A1(Out_Exponent[1]), .A2(n837), .ZN(out[24]) );
  BUF_X1 U664 ( .A(n6), .Z(n138) );
  BUF_X1 U665 ( .A(n6), .Z(n130) );
  BUF_X1 U666 ( .A(n6), .Z(n136) );
  BUF_X1 U667 ( .A(n6), .Z(n140) );
  BUF_X1 U668 ( .A(n6), .Z(n137) );
  BUF_X1 U669 ( .A(n6), .Z(n134) );
  BUF_X1 U670 ( .A(n6), .Z(n135) );
  BUF_X1 U671 ( .A(n6), .Z(n133) );
  BUF_X1 U672 ( .A(n6), .Z(n132) );
  BUF_X1 U673 ( .A(n6), .Z(n131) );
  INV_X1 U674 ( .A(overFlow), .ZN(n837) );
  NOR3_X1 U675 ( .A1(n361), .A2(overFlow), .A3(n362), .ZN(out[31]) );
  NOR4_X1 U676 ( .A1(n363), .A2(n364), .A3(n365), .A4(n366), .ZN(n361) );
  NAND3_X1 U677 ( .A1(n367), .A2(n368), .A3(n369), .ZN(n366) );
  NAND4_X1 U678 ( .A1(n372), .A2(n373), .A3(n374), .A4(n375), .ZN(n364) );
  INV_X1 U679 ( .A(in2[20]), .ZN(n245) );
  INV_X1 U680 ( .A(in2[18]), .ZN(n244) );
  INV_X1 U681 ( .A(in2[16]), .ZN(n243) );
  INV_X1 U682 ( .A(in2[14]), .ZN(n242) );
  INV_X1 U683 ( .A(in2[12]), .ZN(n241) );
  INV_X1 U684 ( .A(in2[10]), .ZN(n240) );
  INV_X1 U685 ( .A(in2[4]), .ZN(n237) );
  INV_X1 U686 ( .A(in2[6]), .ZN(n238) );
  INV_X1 U687 ( .A(in2[8]), .ZN(n239) );
  AOI21_X1 U688 ( .B1(N99), .B2(N97), .A(N31), .ZN(n3530) );
  INV_X1 U689 ( .A(n356), .ZN(sub_64_aco_A_6_) );
  AOI22_X1 U690 ( .A1(n139), .A2(N230), .B1(n128), .B2(N197), .ZN(n356) );
  OR2_X1 U691 ( .A1(N552), .A2(sub_64_I9_aco_carry[1]), .ZN(
        sub_64_I9_aco_carry[2]) );
  OR2_X1 U692 ( .A1(N620), .A2(sub_64_I11_aco_carry[1]), .ZN(
        sub_64_I11_aco_carry[2]) );
  OR2_X1 U693 ( .A1(N688), .A2(sub_64_I13_aco_carry[1]), .ZN(
        sub_64_I13_aco_carry[2]) );
  OR2_X1 U694 ( .A1(N484), .A2(sub_64_I7_aco_carry[1]), .ZN(
        sub_64_I7_aco_carry[2]) );
  OR2_X1 U695 ( .A1(n630), .A2(N313), .ZN(sub_64_I2_aco_carry[1]) );
  OR2_X1 U696 ( .A1(n628), .A2(N381), .ZN(sub_64_I4_aco_carry[1]) );
  OR2_X1 U697 ( .A1(N756), .A2(sub_64_I15_aco_carry[1]), .ZN(
        sub_64_I15_aco_carry[2]) );
  OR2_X1 U698 ( .A1(N416), .A2(sub_64_I5_aco_carry[1]), .ZN(
        sub_64_I5_aco_carry[2]) );
  OR2_X1 U699 ( .A1(n600), .A2(N517), .ZN(sub_64_I8_aco_carry[1]) );
  OR2_X1 U700 ( .A1(N348), .A2(sub_64_I3_aco_carry[1]), .ZN(
        sub_64_I3_aco_carry[2]) );
  OR2_X1 U701 ( .A1(n568), .A2(N585), .ZN(sub_64_I10_aco_carry[1]) );
  OR2_X1 U702 ( .A1(N824), .A2(sub_64_I17_aco_carry[1]), .ZN(
        sub_64_I17_aco_carry[2]) );
  OR2_X1 U703 ( .A1(n549), .A2(N653), .ZN(sub_64_I12_aco_carry[1]) );
  OR2_X1 U704 ( .A1(n529), .A2(N721), .ZN(sub_64_I14_aco_carry[1]) );
  OR2_X1 U705 ( .A1(n562), .A2(N789), .ZN(sub_64_I16_aco_carry[1]) );
  INV_X1 U706 ( .A(n358), .ZN(sub_64_aco_A_2_) );
  NAND2_X1 U707 ( .A1(n359), .A2(n11), .ZN(sub_64_aco_carry[2]) );
  AOI22_X1 U708 ( .A1(n138), .A2(N226), .B1(n128), .B2(N193), .ZN(n358) );
  OAI22_X1 U709 ( .A1(n128), .A2(n8), .B1(n139), .B2(n839), .ZN(N258) );
  OAI22_X1 U710 ( .A1(n128), .A2(n9), .B1(n140), .B2(n838), .ZN(N259) );
  OR2_X1 U711 ( .A1(n457), .A2(N925), .ZN(sub_64_I20_aco_carry[1]) );
  OR2_X1 U712 ( .A1(n559), .A2(N857), .ZN(sub_64_I18_aco_carry[1]) );
  OR2_X1 U713 ( .A1(n474), .A2(N891), .ZN(sub_64_I19_aco_carry[1]) );
  INV_X1 U714 ( .A(n357), .ZN(sub_64_aco_A_5_) );
  AOI22_X1 U715 ( .A1(n139), .A2(N229), .B1(n128), .B2(N196), .ZN(n357) );
  OR2_X1 U716 ( .A1(N960), .A2(sub_64_I21_aco_carry[1]), .ZN(
        sub_64_I21_aco_carry[2]) );
  OR2_X1 U717 ( .A1(n582), .A2(N993), .ZN(sub_64_I22_aco_carry[1]) );
  OR2_X1 U718 ( .A1(n6240), .A2(N449), .ZN(sub_64_I6_aco_carry[1]) );
  AND2_X1 U719 ( .A1(add_42_B_0_), .A2(n84), .ZN(n10) );
  INV_X1 U720 ( .A(in1[2]), .ZN(n2250) );
  INV_X1 U721 ( .A(in1[1]), .ZN(n2240) );
  INV_X1 U722 ( .A(in1[3]), .ZN(n2260) );
  AOI22_X1 U723 ( .A1(n60), .A2(in2[31]), .B1(n33), .B2(in1[31]), .ZN(n362) );
  INV_X1 U724 ( .A(n1800), .ZN(n1940) );
  INV_X1 U725 ( .A(in1[16]), .ZN(n887) );
  INV_X1 U726 ( .A(in1[18]), .ZN(n886) );
  INV_X1 U727 ( .A(in2[13]), .ZN(n868) );
  INV_X1 U728 ( .A(in1[12]), .ZN(n889) );
  INV_X1 U729 ( .A(in1[14]), .ZN(n888) );
  INV_X1 U730 ( .A(in2[15]), .ZN(n867) );
  INV_X1 U731 ( .A(in2[11]), .ZN(n869) );
  INV_X1 U732 ( .A(in1[10]), .ZN(n890) );
  INV_X1 U733 ( .A(in1[0]), .ZN(n8940) );
  AOI22_X1 U734 ( .A1(in2[31]), .A2(n32), .B1(in1[31]), .B2(n142), .ZN(n805)
         );
  INV_X1 U735 ( .A(in2[17]), .ZN(n866) );
  INV_X1 U736 ( .A(in1[6]), .ZN(n8920) );
  INV_X1 U737 ( .A(in1[4]), .ZN(n8930) );
  INV_X1 U738 ( .A(in1[8]), .ZN(n8910) );
  INV_X1 U739 ( .A(in1[20]), .ZN(n884) );
  INV_X1 U740 ( .A(in1[19]), .ZN(n885) );
  INV_X1 U741 ( .A(in2[3]), .ZN(n873) );
  INV_X1 U742 ( .A(in2[19]), .ZN(n865) );
  INV_X1 U743 ( .A(in2[7]), .ZN(n871) );
  INV_X1 U744 ( .A(in2[5]), .ZN(n872) );
  INV_X1 U745 ( .A(in2[21]), .ZN(n8640) );
  INV_X1 U746 ( .A(in1[22]), .ZN(n883) );
  INV_X1 U747 ( .A(in1[27]), .ZN(n878) );
  INV_X1 U748 ( .A(in2[2]), .ZN(n874) );
  INV_X1 U749 ( .A(in2[1]), .ZN(n875) );
  INV_X1 U750 ( .A(in1[24]), .ZN(n881) );
  INV_X1 U751 ( .A(in2[9]), .ZN(n870) );
  INV_X1 U752 ( .A(in1[25]), .ZN(n880) );
  INV_X1 U753 ( .A(in1[26]), .ZN(n879) );
  INV_X1 U754 ( .A(in2[25]), .ZN(n1960) );
  INV_X1 U755 ( .A(in2[27]), .ZN(n1980) );
  INV_X1 U756 ( .A(in2[24]), .ZN(n1950) );
  INV_X1 U757 ( .A(in2[26]), .ZN(n1970) );
  INV_X1 U758 ( .A(in2[28]), .ZN(n199) );
  INV_X1 U759 ( .A(in2[22]), .ZN(n246) );
  INV_X1 U760 ( .A(in1[23]), .ZN(n882) );
  INV_X1 U761 ( .A(in2[23]), .ZN(n1930) );
  INV_X1 U762 ( .A(in1[29]), .ZN(n1920) );
  INV_X1 U763 ( .A(in2[30]), .ZN(n200) );
  INV_X1 U764 ( .A(in1[9]), .ZN(n2290) );
  INV_X1 U765 ( .A(in1[21]), .ZN(n234) );
  INV_X1 U766 ( .A(in1[17]), .ZN(n233) );
  INV_X1 U767 ( .A(in1[15]), .ZN(n232) );
  INV_X1 U768 ( .A(in1[13]), .ZN(n2310) );
  INV_X1 U769 ( .A(in1[11]), .ZN(n2300) );
  INV_X1 U770 ( .A(in1[5]), .ZN(n227) );
  INV_X1 U771 ( .A(in1[7]), .ZN(n228) );
  INV_X1 U772 ( .A(in1[28]), .ZN(n877) );
  INV_X1 U773 ( .A(in2[29]), .ZN(n8630) );
  INV_X1 U774 ( .A(in1[30]), .ZN(n876) );
  AND2_X1 U775 ( .A1(Out_Exponent[6]), .A2(n837), .ZN(out[29]) );
  XOR2_X2 U776 ( .A(n571), .B(n77), .Z(n468) );
  NOR2_X2 U777 ( .A1(n571), .A2(n77), .ZN(n466) );
  CLKBUF_X1 U778 ( .A(n474), .Z(n15) );
  OAI221_X1 U779 ( .B1(n665), .B2(n666), .C1(n295), .C2(n66), .A(n296), .ZN(
        n474) );
  INV_X1 U780 ( .A(n15), .ZN(sub_64_I19_aco_B_0_) );
  INV_X1 U781 ( .A(n511), .ZN(sub_64_I15_aco_B_0_) );
  NAND2_X1 U782 ( .A1(n82), .A2(n530), .ZN(n546) );
  OAI221_X1 U783 ( .B1(n818), .B2(n423), .C1(n528), .C2(n530), .A(n531), .ZN(
        n513) );
  NAND3_X1 U784 ( .A1(n515), .A2(n530), .A3(sub_64_I12_aco_B_0_), .ZN(n531) );
  NAND2_X1 U785 ( .A1(n530), .A2(n76), .ZN(n423) );
  OAI221_X1 U786 ( .B1(n579), .B2(n576), .C1(n608), .C2(n609), .A(n610), .ZN(
        n5560) );
  INV_X1 U787 ( .A(n609), .ZN(sub_64_I3_aco_B_0_) );
  OAI21_X1 U788 ( .B1(sub_64_I3_aco_B_0_), .B2(n608), .A(n629), .ZN(n574) );
  CLKBUF_X1 U789 ( .A(sub_64_I21_aco_B_0_), .Z(n16) );
  CLKBUF_X1 U790 ( .A(sub_64_I21_aco_B_0_), .Z(n17) );
  INV_X1 U791 ( .A(n4550), .ZN(sub_64_I21_aco_B_0_) );
  AOI21_X1 U792 ( .B1(n4900), .B2(n560), .A(n616), .ZN(n5890) );
  OAI221_X1 U793 ( .B1(n324), .B2(n401), .C1(n311), .C2(n4900), .A(n491), .ZN(
        n477) );
  NAND2_X1 U794 ( .A1(n4900), .A2(n78), .ZN(n401) );
  XOR2_X2 U795 ( .A(n4900), .B(sub_64_I16_aco_B_0_), .Z(n403) );
  CLKBUF_X1 U796 ( .A(sub_64_I13_aco_B_0_), .Z(n18) );
  CLKBUF_X1 U797 ( .A(sub_64_I13_aco_B_0_), .Z(n19) );
  INV_X1 U798 ( .A(n530), .ZN(sub_64_I13_aco_B_0_) );
  OAI22_X1 U799 ( .A1(n44), .A2(n233), .B1(n56), .B2(n866), .ZN(inShift[17])
         );
  CLKBUF_X1 U800 ( .A(n3530), .Z(n20) );
  INV_X1 U801 ( .A(n22), .ZN(n60) );
  OAI22_X1 U802 ( .A1(n22), .A2(n1930), .B1(n58), .B2(n882), .ZN(a[23]) );
  INV_X1 U803 ( .A(b[24]), .ZN(n148) );
  BUF_X1 U804 ( .A(n3530), .Z(n22) );
  CLKBUF_X1 U805 ( .A(a[23]), .Z(n84) );
  INV_X1 U806 ( .A(n60), .ZN(n23) );
  INV_X1 U807 ( .A(n59), .ZN(n24) );
  INV_X1 U808 ( .A(n60), .ZN(n25) );
  INV_X1 U809 ( .A(n56), .ZN(n26) );
  INV_X1 U810 ( .A(n65), .ZN(n27) );
  INV_X1 U811 ( .A(n65), .ZN(n28) );
  INV_X1 U812 ( .A(n65), .ZN(n29) );
  INV_X1 U813 ( .A(n65), .ZN(n30) );
  INV_X1 U814 ( .A(n64), .ZN(n3100) );
  INV_X1 U815 ( .A(n64), .ZN(n32) );
  INV_X1 U816 ( .A(n64), .ZN(n33) );
  INV_X1 U817 ( .A(n64), .ZN(n34) );
  INV_X1 U818 ( .A(n61), .ZN(n35) );
  INV_X1 U819 ( .A(n60), .ZN(n36) );
  INV_X1 U820 ( .A(n61), .ZN(n37) );
  INV_X1 U821 ( .A(n143), .ZN(n38) );
  INV_X1 U822 ( .A(n144), .ZN(n39) );
  INV_X1 U823 ( .A(n144), .ZN(n40) );
  INV_X1 U824 ( .A(n144), .ZN(n41) );
  INV_X1 U825 ( .A(n142), .ZN(n42) );
  INV_X1 U826 ( .A(n142), .ZN(n43) );
  INV_X1 U827 ( .A(n142), .ZN(n44) );
  INV_X1 U828 ( .A(n142), .ZN(n45) );
  INV_X1 U829 ( .A(n145), .ZN(n46) );
  INV_X1 U830 ( .A(n145), .ZN(n47) );
  INV_X1 U831 ( .A(n145), .ZN(n48) );
  INV_X1 U832 ( .A(n145), .ZN(n49) );
  INV_X1 U833 ( .A(n61), .ZN(n50) );
  INV_X1 U834 ( .A(n60), .ZN(n51) );
  INV_X1 U835 ( .A(n61), .ZN(n52) );
  INV_X1 U836 ( .A(n60), .ZN(n53) );
  INV_X1 U837 ( .A(n24), .ZN(n54) );
  INV_X1 U838 ( .A(n141), .ZN(n55) );
  INV_X1 U839 ( .A(n21), .ZN(n56) );
  INV_X1 U840 ( .A(n21), .ZN(n57) );
  INV_X1 U841 ( .A(n3530), .ZN(n58) );
  INV_X1 U842 ( .A(n21), .ZN(n59) );
  INV_X1 U843 ( .A(n22), .ZN(n61) );
  CLKBUF_X1 U844 ( .A(n59), .Z(n65) );
  CLKBUF_X1 U845 ( .A(n59), .Z(n64) );
  INV_X1 U846 ( .A(n146), .ZN(n145) );
  NAND4_X1 U847 ( .A1(n8), .A2(n9), .A3(n802), .A4(n803), .ZN(n798) );
  INV_X1 U848 ( .A(n568), .ZN(sub_64_I10_aco_B_0_) );
  NAND2_X1 U849 ( .A1(n18), .A2(sub_64_I12_aco_B_0_), .ZN(n424) );
  OR4_X1 U850 ( .A1(N658), .A2(N657), .A3(N660), .A4(N659), .ZN(n733) );
  NAND3_X1 U851 ( .A1(n16), .A2(n583), .A3(n249), .ZN(n5850) );
  NAND2_X1 U852 ( .A1(n248), .A2(n16), .ZN(n4520) );
  NOR3_X1 U853 ( .A1(n411), .A2(n18), .A3(n595), .ZN(n615) );
  INV_X1 U854 ( .A(n76), .ZN(sub_64_I12_aco_B_0_) );
  INV_X1 U855 ( .A(n630), .ZN(sub_64_I2_aco_B_0_) );
  NOR3_X1 U856 ( .A1(n286), .A2(n17), .A3(n80), .ZN(n4560) );
  AOI22_X1 U862 ( .A1(n83), .A2(n598), .B1(sub_64_I10_aco_B_0_), .B2(n8270), 
        .ZN(n597) );
  AOI22_X1 U863 ( .A1(n598), .A2(sub_64_I10_aco_B_0_), .B1(n83), .B2(n569), 
        .ZN(n567) );
  AOI22_X1 U864 ( .A1(n83), .A2(n8260), .B1(n569), .B2(sub_64_I10_aco_B_0_), 
        .ZN(n5510) );
  NAND3_X1 U865 ( .A1(n473), .A2(n15), .A3(sub_64_I20_aco_B_0_), .ZN(n472) );
  NAND2_X1 U866 ( .A1(n16), .A2(sub_64_I20_aco_B_0_), .ZN(n3880) );
  OR4_X1 U867 ( .A1(N862), .A2(N861), .A3(N864), .A4(N863), .ZN(n667) );
  OAI21_X1 U868 ( .B1(n636), .B2(n637), .A(n250), .ZN(n582) );
  CLKBUF_X1 U869 ( .A(sub_64_I18_aco_B_0_), .Z(n62) );
  CLKBUF_X1 U870 ( .A(sub_64_I18_aco_B_0_), .Z(n63) );
  INV_X1 U871 ( .A(n559), .ZN(sub_64_I18_aco_B_0_) );
  INV_X1 U872 ( .A(n146), .ZN(n144) );
  CLKBUF_X1 U873 ( .A(n559), .Z(n66) );
  OAI21_X1 U874 ( .B1(n667), .B2(n668), .A(n296), .ZN(n559) );
  INV_X1 U875 ( .A(n606), .ZN(sub_64_I5_aco_B_0_) );
  OR3_X1 U876 ( .A1(n528), .A2(n18), .A3(n82), .ZN(n527) );
  INV_X1 U877 ( .A(n582), .ZN(sub_64_I22_aco_B_0_) );
  OR4_X1 U878 ( .A1(N522), .A2(N521), .A3(N524), .A4(N523), .ZN(n764) );
  CLKBUF_X1 U879 ( .A(sub_64_I9_aco_B_0_), .Z(n67) );
  INV_X1 U880 ( .A(n571), .ZN(sub_64_I9_aco_B_0_) );
  INV_X1 U881 ( .A(n5520), .ZN(sub_64_I11_aco_B_0_) );
  NAND2_X1 U882 ( .A1(n5520), .A2(n83), .ZN(n438) );
  NAND3_X1 U883 ( .A1(n8260), .A2(n5520), .A3(sub_64_I10_aco_B_0_), .ZN(n5530)
         );
  OAI221_X1 U884 ( .B1(n5170), .B2(n124), .C1(n5510), .C2(n5520), .A(n5530), 
        .ZN(n515) );
  NAND3_X1 U885 ( .A1(n835), .A2(n609), .A3(sub_64_I2_aco_B_0_), .ZN(n610) );
  NAND2_X1 U886 ( .A1(sub_64_I3_aco_B_0_), .A2(sub_64_I2_aco_B_0_), .ZN(n91)
         );
  NAND2_X1 U887 ( .A1(sub_64_I3_aco_B_0_), .A2(sub_64_I2_aco_B_0_), .ZN(n578)
         );
  INV_X1 U888 ( .A(n6240), .ZN(sub_64_I6_aco_B_0_) );
  NAND2_X1 U889 ( .A1(sub_64_I7_aco_B_0_), .A2(sub_64_I6_aco_B_0_), .ZN(n108)
         );
  NAND2_X1 U890 ( .A1(sub_64_I7_aco_B_0_), .A2(sub_64_I6_aco_B_0_), .ZN(n109)
         );
  NAND2_X1 U891 ( .A1(sub_64_I7_aco_B_0_), .A2(sub_64_I6_aco_B_0_), .ZN(n501)
         );
  NOR2_X1 U892 ( .A1(n6230), .A2(sub_64_I7_aco_B_0_), .ZN(n6220) );
  INV_X1 U893 ( .A(n603), .ZN(sub_64_I7_aco_B_0_) );
  OR4_X1 U894 ( .A1(N828), .A2(N827), .A3(N830), .A4(N829), .ZN(n6880) );
  INV_X1 U895 ( .A(sub_64_aco_B_0_), .ZN(n68) );
  INV_X1 U896 ( .A(n68), .ZN(n69) );
  INV_X1 U897 ( .A(n68), .ZN(n70) );
  INV_X1 U898 ( .A(n68), .ZN(n71) );
  INV_X1 U899 ( .A(n126), .ZN(n72) );
  INV_X1 U900 ( .A(n72), .ZN(n73) );
  INV_X1 U901 ( .A(n72), .ZN(n74) );
  INV_X1 U902 ( .A(n72), .ZN(n75) );
  INV_X1 U903 ( .A(n127), .ZN(n126) );
  OR3_X1 U904 ( .A1(n3870), .A2(sub_64_I19_aco_B_0_), .A3(n5870), .ZN(n611) );
  NAND2_X1 U905 ( .A1(sub_64_I20_aco_B_0_), .A2(sub_64_I19_aco_B_0_), .ZN(n471) );
  OAI21_X1 U906 ( .B1(sub_46_ni_B_0_), .B2(n371), .A(n635), .ZN(n632) );
  NAND3_X1 U907 ( .A1(n128), .A2(sub_46_ni_B_0_), .A3(N165), .ZN(n635) );
  NAND2_X1 U908 ( .A1(N188), .A2(n129), .ZN(sub_46_ni_B_0_) );
  CLKBUF_X1 U909 ( .A(n549), .Z(n76) );
  OAI21_X1 U910 ( .B1(n733), .B2(n734), .A(n809), .ZN(n549) );
  AOI21_X1 U911 ( .B1(n6240), .B2(n573), .A(n6250), .ZN(n602) );
  NAND3_X1 U912 ( .A1(n990), .A2(n6240), .A3(n6260), .ZN(n6230) );
  NAND2_X1 U913 ( .A1(sub_64_I17_aco_B_0_), .A2(sub_64_I16_aco_B_0_), .ZN(n402) );
  CLKBUF_X1 U914 ( .A(n600), .Z(n77) );
  OAI21_X1 U915 ( .B1(n764), .B2(n765), .A(n8300), .ZN(n600) );
  NAND2_X1 U916 ( .A1(n609), .A2(n630), .ZN(n576) );
  NAND2_X1 U917 ( .A1(n609), .A2(n630), .ZN(n90) );
  NAND3_X1 U918 ( .A1(sub_64_I3_aco_B_0_), .A2(n630), .A3(n836), .ZN(n629) );
  AOI22_X1 U919 ( .A1(n630), .A2(n835), .B1(sub_64_I2_aco_B_0_), .B2(n836), 
        .ZN(n608) );
  NOR2_X1 U920 ( .A1(n606), .A2(n628), .ZN(n539) );
  AND3_X1 U921 ( .A1(n574), .A2(n606), .A3(sub_64_I4_aco_B_0_), .ZN(n605) );
  CLKBUF_X1 U922 ( .A(n562), .Z(n78) );
  OAI21_X1 U923 ( .B1(n6900), .B2(n6910), .A(n3190), .ZN(n562) );
  CLKBUF_X1 U924 ( .A(n457), .Z(n80) );
  OAI21_X1 U925 ( .B1(n641), .B2(n642), .A(n274), .ZN(n457) );
  CLKBUF_X1 U926 ( .A(n529), .Z(n82) );
  OAI21_X1 U927 ( .B1(n713), .B2(n714), .A(n342), .ZN(n529) );
  CLKBUF_X1 U928 ( .A(n568), .Z(n83) );
  OAI21_X1 U929 ( .B1(n751), .B2(n752), .A(n738), .ZN(n568) );
  INV_X1 U930 ( .A(n628), .ZN(sub_64_I4_aco_B_0_) );
  OAI21_X1 U931 ( .B1(n787), .B2(n788), .A(n834), .ZN(n628) );
  INV_X1 U932 ( .A(n2030), .ZN(n236) );
  AND2_X1 U933 ( .A1(Out_Exponent[7]), .A2(n837), .ZN(out[30]) );
  NAND2_X1 U934 ( .A1(n632), .A2(n127), .ZN(n631) );
  NAND4_X1 U935 ( .A1(n370), .A2(n798), .A3(n799), .A4(sub_46_ni_B_0_), .ZN(
        n634) );
  OAI22_X1 U936 ( .A1(n38), .A2(n870), .B1(n143), .B2(n2290), .ZN(a[9]) );
  OAI22_X1 U937 ( .A1(n38), .A2(n239), .B1(n54), .B2(n8910), .ZN(a[8]) );
  OAI22_X1 U938 ( .A1(n38), .A2(n871), .B1(n55), .B2(n228), .ZN(a[7]) );
  OAI22_X1 U939 ( .A1(n38), .A2(n238), .B1(n56), .B2(n8920), .ZN(a[6]) );
  OAI22_X1 U940 ( .A1(n38), .A2(n872), .B1(n57), .B2(n227), .ZN(a[5]) );
  OAI22_X1 U941 ( .A1(n38), .A2(n237), .B1(n58), .B2(n8930), .ZN(a[4]) );
  OAI22_X1 U942 ( .A1(n39), .A2(n873), .B1(n143), .B2(n2260), .ZN(a[3]) );
  OAI22_X1 U943 ( .A1(n50), .A2(n2290), .B1(n55), .B2(n870), .ZN(inShift[9])
         );
  OAI22_X1 U944 ( .A1(n46), .A2(n879), .B1(n142), .B2(n1970), .ZN(b[26]) );
  OAI22_X1 U945 ( .A1(n141), .A2(n880), .B1(n59), .B2(n1960), .ZN(b[25]) );
  OAI22_X1 U946 ( .A1(n26), .A2(n881), .B1(n57), .B2(n1950), .ZN(b[24]) );
  OR4_X1 U947 ( .A1(N420), .A2(N419), .A3(N422), .A4(N421), .ZN(n785) );
  AND3_X1 U948 ( .A1(n5540), .A2(n571), .A3(sub_64_I8_aco_B_0_), .ZN(n570) );
  OAI22_X1 U949 ( .A1(n67), .A2(n572), .B1(n599), .B2(n571), .ZN(n569) );
  NAND2_X1 U950 ( .A1(sub_64_I14_aco_B_0_), .A2(n19), .ZN(n526) );
  OAI221_X1 U951 ( .B1(n525), .B2(n526), .C1(sub_64_I14_aco_B_0_), .C2(n806), 
        .A(n527), .ZN(n510) );
  INV_X1 U952 ( .A(n82), .ZN(sub_64_I14_aco_B_0_) );
  OR4_X1 U953 ( .A1(N896), .A2(N895), .A3(N898), .A4(N897), .ZN(n665) );
  INV_X1 U954 ( .A(in2[0]), .ZN(n235) );
  OR4_X1 U955 ( .A1(N556), .A2(N555), .A3(N558), .A4(N557), .ZN(n7620) );
  INV_X1 U956 ( .A(sub_64_aco_B_0_), .ZN(n127) );
  INV_X1 U957 ( .A(n634), .ZN(sub_64_aco_B_0_) );
  OAI22_X1 U958 ( .A1(n30), .A2(n8630), .B1(n54), .B2(n1920), .ZN(a[29]) );
  OAI22_X1 U959 ( .A1(n49), .A2(n199), .B1(n55), .B2(n877), .ZN(a[28]) );
  OAI22_X1 U960 ( .A1(n50), .A2(n246), .B1(n56), .B2(n883), .ZN(a[22]) );
  OAI22_X1 U961 ( .A1(n51), .A2(n8640), .B1(n57), .B2(n234), .ZN(a[21]) );
  OAI22_X1 U962 ( .A1(n3100), .A2(n245), .B1(n58), .B2(n884), .ZN(a[20]) );
  OAI22_X1 U963 ( .A1(n52), .A2(n865), .B1(n143), .B2(n885), .ZN(a[19]) );
  OAI22_X1 U964 ( .A1(n40), .A2(n874), .B1(n142), .B2(n2250), .ZN(a[2]) );
  OAI22_X1 U965 ( .A1(n41), .A2(n875), .B1(n143), .B2(n2240), .ZN(a[1]) );
  OAI22_X1 U966 ( .A1(n29), .A2(n1980), .B1(n143), .B2(n878), .ZN(a[27]) );
  OAI22_X1 U967 ( .A1(n24), .A2(n1970), .B1(n58), .B2(n879), .ZN(a[26]) );
  OAI22_X1 U968 ( .A1(n146), .A2(n1960), .B1(n55), .B2(n880), .ZN(a[25]) );
  OAI22_X1 U969 ( .A1(n21), .A2(n1950), .B1(n56), .B2(n881), .ZN(a[24]) );
  OAI22_X1 U970 ( .A1(n22), .A2(n882), .B1(n58), .B2(n1930), .ZN(b[23]) );
  INV_X1 U971 ( .A(b[23]), .ZN(n147) );
  OAI221_X4 U972 ( .B1(n774), .B2(n775), .C1(n767), .C2(n6240), .A(n768), .ZN(
        n603) );
  NAND3_X1 U973 ( .A1(n4540), .A2(n4550), .A3(n248), .ZN(n4530) );
  AOI21_X1 U974 ( .B1(n4550), .B2(n583), .A(n612), .ZN(n584) );
  NAND2_X1 U975 ( .A1(n249), .A2(n4550), .ZN(n470) );
  NOR3_X1 U976 ( .A1(n4850), .A2(n4550), .A3(n5870), .ZN(n612) );
  NAND2_X1 U977 ( .A1(n4550), .A2(n80), .ZN(n3870) );
  AOI21_X1 U978 ( .B1(n511), .B2(n563), .A(n617), .ZN(n5920) );
  NOR3_X1 U979 ( .A1(n546), .A2(n511), .A3(n595), .ZN(n617) );
  NAND2_X1 U980 ( .A1(n78), .A2(n511), .ZN(n5230) );
  OAI221_X1 U981 ( .B1(n3490), .B2(n411), .C1(n335), .C2(n511), .A(n512), .ZN(
        n492) );
  NAND3_X1 U982 ( .A1(n513), .A2(n511), .A3(sub_64_I14_aco_B_0_), .ZN(n512) );
  OAI22_X1 U983 ( .A1(sub_64_I11_aco_B_0_), .A2(n567), .B1(n597), .B2(n5520), 
        .ZN(n566) );
  AOI22_X1 U984 ( .A1(n77), .A2(n601), .B1(sub_64_I8_aco_B_0_), .B2(n6220), 
        .ZN(n599) );
  AOI22_X1 U985 ( .A1(n77), .A2(n5540), .B1(n601), .B2(sub_64_I8_aco_B_0_), 
        .ZN(n572) );
  OAI22_X1 U986 ( .A1(sub_64_I7_aco_B_0_), .A2(n602), .B1(n603), .B2(n6230), 
        .ZN(n601) );
  OAI221_X1 U987 ( .B1(n5550), .B2(n499), .C1(n602), .C2(n603), .A(n604), .ZN(
        n5540) );
  NAND3_X1 U988 ( .A1(n573), .A2(n603), .A3(sub_64_I6_aco_B_0_), .ZN(n604) );
  NAND2_X1 U989 ( .A1(n603), .A2(n6240), .ZN(n107) );
  NAND2_X1 U990 ( .A1(n603), .A2(n6240), .ZN(n499) );
  OAI22_X1 U991 ( .A1(n27), .A2(n200), .B1(n143), .B2(n876), .ZN(a[30]) );
  INV_X1 U992 ( .A(n223), .ZN(n247) );
  OR4_X1 U993 ( .A1(N760), .A2(N759), .A3(N762), .A4(N761), .ZN(n711) );
  OR4_X1 U994 ( .A1(N488), .A2(N487), .A3(N490), .A4(N489), .ZN(n774) );
  OR4_X1 U995 ( .A1(N624), .A2(N623), .A3(N626), .A4(N625), .ZN(n749) );
  OR4_X1 U996 ( .A1(N964), .A2(N963), .A3(N966), .A4(N965), .ZN(n639) );
  OR4_X1 U997 ( .A1(N454), .A2(N453), .A3(N456), .A4(N455), .ZN(n776) );
  OR4_X1 U998 ( .A1(N794), .A2(N793), .A3(N796), .A4(N795), .ZN(n6900) );
  OR4_X1 U999 ( .A1(N386), .A2(N385), .A3(N388), .A4(N387), .ZN(n787) );
  OR4_X1 U1000 ( .A1(N692), .A2(N691), .A3(N694), .A4(N693), .ZN(n731) );
  OR4_X1 U1001 ( .A1(N930), .A2(N929), .A3(N932), .A4(N931), .ZN(n641) );
  OR4_X1 U1002 ( .A1(N590), .A2(N589), .A3(N592), .A4(N591), .ZN(n751) );
  OR4_X1 U1003 ( .A1(N726), .A2(N725), .A3(N728), .A4(N727), .ZN(n713) );
  OR4_X1 U1004 ( .A1(N352), .A2(N351), .A3(N354), .A4(N353), .ZN(n7940) );
  INV_X1 U1005 ( .A(n4900), .ZN(sub_64_I17_aco_B_0_) );
  INV_X1 U1006 ( .A(n80), .ZN(sub_64_I20_aco_B_0_) );
  INV_X1 U1007 ( .A(n78), .ZN(sub_64_I16_aco_B_0_) );
  INV_X1 U1008 ( .A(sub_46_ni_B_0_), .ZN(add_42_B_0_) );
  OR4_X1 U1009 ( .A1(N318), .A2(N317), .A3(N320), .A4(N319), .ZN(n7960) );
  OR4_X1 U1010 ( .A1(N993), .A2(N1000), .A3(N995), .A4(N994), .ZN(n637) );
  NOR3_X1 U1011 ( .A1(N196), .A2(N198), .A3(N197), .ZN(n800) );
  NAND4_X1 U1012 ( .A1(n839), .A2(n838), .A3(n800), .A4(n801), .ZN(n799) );
  NAND3_X1 U1013 ( .A1(n309), .A2(n66), .A3(n615), .ZN(n5870) );
  OAI21_X1 U1014 ( .B1(n62), .B2(n5890), .A(n614), .ZN(n613) );
  OAI221_X1 U1015 ( .B1(n3160), .B2(n506), .C1(n5890), .C2(n66), .A(n5900), 
        .ZN(n5880) );
  NAND3_X1 U1016 ( .A1(n63), .A2(n309), .A3(n615), .ZN(n614) );
  NAND3_X1 U1017 ( .A1(n560), .A2(n66), .A3(sub_64_I17_aco_B_0_), .ZN(n5900)
         );
  NAND3_X1 U1018 ( .A1(n477), .A2(n15), .A3(n62), .ZN(n476) );
  NAND2_X1 U1019 ( .A1(n66), .A2(n4900), .ZN(n506) );
  NOR3_X1 U1020 ( .A1(n4900), .A2(sub_64_I16_aco_B_0_), .A3(n333), .ZN(n616)
         );
  OAI22_X1 U1021 ( .A1(sub_64_I16_aco_B_0_), .A2(n5920), .B1(n78), .B2(n333), 
        .ZN(n560) );
  NAND3_X1 U1022 ( .A1(n563), .A2(n78), .A3(sub_64_I15_aco_B_0_), .ZN(n593) );
  NAND3_X1 U1023 ( .A1(n4890), .A2(n4900), .A3(n63), .ZN(n4880) );
  NAND2_X1 U1024 ( .A1(n62), .A2(sub_64_I17_aco_B_0_), .ZN(n4870) );
  NAND3_X1 U1025 ( .A1(n492), .A2(n4900), .A3(sub_64_I16_aco_B_0_), .ZN(n491)
         );
  NAND3_X1 U1026 ( .A1(n510), .A2(n511), .A3(sub_64_I16_aco_B_0_), .ZN(n509)
         );
  NAND2_X1 U1027 ( .A1(sub_64_I16_aco_B_0_), .A2(sub_64_I15_aco_B_0_), .ZN(
        n508) );
  NAND2_X1 U1028 ( .A1(n15), .A2(n66), .ZN(n393) );
  NAND2_X1 U1029 ( .A1(sub_64_I19_aco_B_0_), .A2(n62), .ZN(n394) );
  NAND2_X1 U1030 ( .A1(sub_64_I15_aco_B_0_), .A2(sub_64_I14_aco_B_0_), .ZN(
        n412) );
  XOR2_X1 U1031 ( .A(n609), .B(sub_64_I2_aco_B_0_), .Z(n85) );
  XOR2_X2 U1032 ( .A(n5520), .B(sub_64_I10_aco_B_0_), .Z(n442) );
  XOR2_X2 U1033 ( .A(n76), .B(n19), .Z(n425) );
  XOR2_X2 U1034 ( .A(n82), .B(sub_64_I15_aco_B_0_), .Z(n413) );
  BUF_X1 U1035 ( .A(n92), .Z(n94) );
  BUF_X1 U1036 ( .A(n92), .Z(n95) );
  BUF_X1 U1037 ( .A(n92), .Z(n96) );
  BUF_X1 U1038 ( .A(n92), .Z(n970) );
  BUF_X1 U1039 ( .A(n93), .Z(n98) );
  BUF_X1 U1040 ( .A(n93), .Z(n990) );
  BUF_X1 U1041 ( .A(n93), .Z(n100) );
  BUF_X1 U1042 ( .A(n93), .Z(n101) );
  BUF_X1 U1043 ( .A(n537), .Z(n102) );
  BUF_X1 U1044 ( .A(n537), .Z(n103) );
  INV_X1 U1045 ( .A(n110), .ZN(n111) );
  INV_X1 U1046 ( .A(n110), .ZN(n112) );
  INV_X1 U1047 ( .A(n111), .ZN(n113) );
  INV_X1 U1048 ( .A(n112), .ZN(n114) );
  INV_X1 U1049 ( .A(n112), .ZN(n115) );
  INV_X1 U1050 ( .A(n464), .ZN(n116) );
  INV_X1 U1051 ( .A(n464), .ZN(n117) );
  INV_X1 U1052 ( .A(n116), .ZN(n118) );
  INV_X1 U1053 ( .A(n116), .ZN(n119) );
  INV_X1 U1054 ( .A(n116), .ZN(n120) );
  INV_X1 U1055 ( .A(n117), .ZN(n121) );
  INV_X1 U1056 ( .A(n146), .ZN(n142) );
  AND2_X1 U1086 ( .A1(in1[23]), .A2(n1930), .ZN(n1740) );
  OAI22_X1 U1087 ( .A1(in1[24]), .A2(n1740), .B1(n1740), .B2(n1950), .ZN(n1750) );
  OR2_X1 U1088 ( .A1(n1920), .A2(in2[29]), .ZN(n1760) );
  NAND2_X1 U1089 ( .A1(in1[28]), .A2(n199), .ZN(n1770) );
  NAND2_X1 U1090 ( .A1(in1[27]), .A2(n1980), .ZN(n1840) );
  NAND4_X1 U1091 ( .A1(n1750), .A2(n1760), .A3(n1770), .A4(n1840), .ZN(n191)
         );
  NAND2_X1 U1092 ( .A1(in1[26]), .A2(n1970), .ZN(n1830) );
  NAND2_X1 U1093 ( .A1(in1[25]), .A2(n1960), .ZN(n1780) );
  NAND2_X1 U1094 ( .A1(n1830), .A2(n1780), .ZN(n190) );
  AND2_X1 U1095 ( .A1(in1[30]), .A2(n200), .ZN(n189) );
  AND2_X1 U1096 ( .A1(n1770), .A2(n1760), .ZN(n1870) );
  NOR2_X1 U1097 ( .A1(n1930), .A2(in1[23]), .ZN(n1800) );
  OAI21_X1 U1098 ( .B1(in1[24]), .B2(n1940), .A(n1950), .ZN(n1790) );
  OAI211_X1 U1099 ( .C1(n1800), .C2(n881), .A(n1790), .B(n1780), .ZN(n1810) );
  OAI221_X1 U1100 ( .B1(in1[25]), .B2(n1960), .C1(in1[26]), .C2(n1970), .A(
        n1810), .ZN(n1820) );
  NAND3_X1 U1101 ( .A1(n1840), .A2(n1830), .A3(n1820), .ZN(n1850) );
  OAI221_X1 U1102 ( .B1(in1[27]), .B2(n1980), .C1(in1[28]), .C2(n199), .A(
        n1850), .ZN(n1860) );
  AOI22_X1 U1103 ( .A1(in2[29]), .A2(n1920), .B1(n1870), .B2(n1860), .ZN(n1880) );
  OAI22_X1 U1104 ( .A1(in1[30]), .A2(n200), .B1(n189), .B2(n1880), .ZN(N31) );
  NOR4_X1 U1105 ( .A1(n191), .A2(n190), .A3(N31), .A4(n189), .ZN(N97) );
  NOR2_X1 U1106 ( .A1(n235), .A2(in1[0]), .ZN(n2020) );
  AND2_X1 U1107 ( .A1(n2240), .A2(n2020), .ZN(n2010) );
  OAI222_X1 U1108 ( .A1(n2020), .A2(n2240), .B1(in2[1]), .B2(n2010), .C1(
        in2[2]), .C2(n2250), .ZN(n2030) );
  AOI221_X1 U1109 ( .B1(n2250), .B2(in2[2]), .C1(n2260), .C2(in2[3]), .A(n236), 
        .ZN(n2040) );
  AOI221_X1 U1110 ( .B1(n873), .B2(in1[3]), .C1(n237), .C2(in1[4]), .A(n2040), 
        .ZN(n2050) );
  AOI221_X1 U1111 ( .B1(n8930), .B2(in2[4]), .C1(n227), .C2(in2[5]), .A(n2050), 
        .ZN(n2060) );
  AOI221_X1 U1112 ( .B1(n872), .B2(in1[5]), .C1(n238), .C2(in1[6]), .A(n2060), 
        .ZN(n2070) );
  AOI221_X1 U1113 ( .B1(n8920), .B2(in2[6]), .C1(n228), .C2(in2[7]), .A(n2070), 
        .ZN(n2080) );
  AOI221_X1 U1114 ( .B1(n871), .B2(in1[7]), .C1(n239), .C2(in1[8]), .A(n2080), 
        .ZN(n2090) );
  AOI221_X1 U1115 ( .B1(n8910), .B2(in2[8]), .C1(n2290), .C2(in2[9]), .A(n2090), .ZN(n2100) );
  AOI221_X1 U1116 ( .B1(n240), .B2(in1[10]), .C1(n870), .C2(in1[9]), .A(n2100), 
        .ZN(n2110) );
  AOI221_X1 U1117 ( .B1(n890), .B2(in2[10]), .C1(n2300), .C2(in2[11]), .A(
        n2110), .ZN(n2120) );
  AOI221_X1 U1118 ( .B1(n869), .B2(in1[11]), .C1(n241), .C2(in1[12]), .A(n2120), .ZN(n2130) );
  AOI221_X1 U1119 ( .B1(n889), .B2(in2[12]), .C1(n2310), .C2(in2[13]), .A(
        n2130), .ZN(n2140) );
  AOI221_X1 U1120 ( .B1(n868), .B2(in1[13]), .C1(n242), .C2(in1[14]), .A(n2140), .ZN(n2150) );
  AOI221_X1 U1121 ( .B1(n888), .B2(in2[14]), .C1(n232), .C2(in2[15]), .A(n2150), .ZN(n2160) );
  AOI221_X1 U1122 ( .B1(n867), .B2(in1[15]), .C1(n243), .C2(in1[16]), .A(n2160), .ZN(n2170) );
  AOI221_X1 U1123 ( .B1(n887), .B2(in2[16]), .C1(n233), .C2(in2[17]), .A(n2170), .ZN(n2180) );
  AOI221_X1 U1124 ( .B1(n866), .B2(in1[17]), .C1(n244), .C2(in1[18]), .A(n2180), .ZN(n2190) );
  AOI221_X1 U1125 ( .B1(n886), .B2(in2[18]), .C1(n885), .C2(in2[19]), .A(n2190), .ZN(n2200) );
  AOI221_X1 U1126 ( .B1(n865), .B2(in1[19]), .C1(n245), .C2(in1[20]), .A(n2200), .ZN(n2210) );
  AOI221_X1 U1127 ( .B1(n884), .B2(in2[20]), .C1(n234), .C2(in2[21]), .A(n2210), .ZN(n2220) );
  AOI221_X1 U1128 ( .B1(n8640), .B2(in1[21]), .C1(n246), .C2(in1[22]), .A(
        n2220), .ZN(n223) );
  OAI21_X1 U1129 ( .B1(in1[22]), .B2(n246), .A(n247), .ZN(N99) );
endmodule


module Register32bit ( clk, rst, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, rst;
  wire   n1;

  DFFR_X1 out_reg_31_ ( .D(in[31]), .CK(clk), .RN(n1), .Q(out[31]) );
  DFFR_X1 out_reg_23_ ( .D(in[23]), .CK(clk), .RN(n1), .Q(out[23]) );
  DFFR_X1 out_reg_0_ ( .D(in[0]), .CK(clk), .RN(n1), .Q(out[0]) );
  DFFR_X1 out_reg_24_ ( .D(in[24]), .CK(clk), .RN(n1), .Q(out[24]) );
  DFFR_X1 out_reg_1_ ( .D(in[1]), .CK(clk), .RN(n1), .Q(out[1]) );
  DFFR_X1 out_reg_22_ ( .D(in[22]), .CK(clk), .RN(n1), .Q(out[22]) );
  DFFR_X1 out_reg_21_ ( .D(in[21]), .CK(clk), .RN(n1), .Q(out[21]) );
  DFFR_X1 out_reg_20_ ( .D(in[20]), .CK(clk), .RN(n1), .Q(out[20]) );
  DFFR_X1 out_reg_19_ ( .D(in[19]), .CK(clk), .RN(n1), .Q(out[19]) );
  DFFR_X1 out_reg_18_ ( .D(in[18]), .CK(clk), .RN(n1), .Q(out[18]) );
  DFFR_X1 out_reg_17_ ( .D(in[17]), .CK(clk), .RN(n1), .Q(out[17]) );
  DFFR_X1 out_reg_16_ ( .D(in[16]), .CK(clk), .RN(n1), .Q(out[16]) );
  DFFR_X1 out_reg_15_ ( .D(in[15]), .CK(clk), .RN(n1), .Q(out[15]) );
  DFFR_X1 out_reg_14_ ( .D(in[14]), .CK(clk), .RN(n1), .Q(out[14]) );
  DFFR_X1 out_reg_13_ ( .D(in[13]), .CK(clk), .RN(n1), .Q(out[13]) );
  DFFR_X1 out_reg_12_ ( .D(in[12]), .CK(clk), .RN(n1), .Q(out[12]) );
  DFFR_X1 out_reg_11_ ( .D(in[11]), .CK(clk), .RN(n1), .Q(out[11]) );
  DFFR_X1 out_reg_10_ ( .D(in[10]), .CK(clk), .RN(n1), .Q(out[10]) );
  DFFR_X1 out_reg_25_ ( .D(in[25]), .CK(clk), .RN(n1), .Q(out[25]) );
  DFFR_X1 out_reg_2_ ( .D(in[2]), .CK(clk), .RN(n1), .Q(out[2]) );
  DFFR_X1 out_reg_8_ ( .D(in[8]), .CK(clk), .RN(n1), .Q(out[8]) );
  DFFR_X1 out_reg_7_ ( .D(in[7]), .CK(clk), .RN(n1), .Q(out[7]) );
  DFFR_X1 out_reg_6_ ( .D(in[6]), .CK(clk), .RN(n1), .Q(out[6]) );
  DFFR_X1 out_reg_5_ ( .D(in[5]), .CK(clk), .RN(n1), .Q(out[5]) );
  DFFR_X1 out_reg_4_ ( .D(in[4]), .CK(clk), .RN(n1), .Q(out[4]) );
  DFFR_X1 out_reg_3_ ( .D(in[3]), .CK(clk), .RN(n1), .Q(out[3]) );
  DFFR_X1 out_reg_9_ ( .D(in[9]), .CK(clk), .RN(n1), .Q(out[9]) );
  DFFR_X1 out_reg_26_ ( .D(in[26]), .CK(clk), .RN(n1), .Q(out[26]) );
  DFFR_X1 out_reg_27_ ( .D(in[27]), .CK(clk), .RN(n1), .Q(out[27]) );
  DFFR_X1 out_reg_28_ ( .D(in[28]), .CK(clk), .RN(n1), .Q(out[28]) );
  DFFR_X1 out_reg_29_ ( .D(in[29]), .CK(clk), .RN(n1), .Q(out[29]) );
  DFFR_X1 out_reg_30_ ( .D(in[30]), .CK(clk), .RN(n1), .Q(out[30]) );
  INV_X2 U3 ( .A(rst), .ZN(n1) );
endmodule


module sync_fpu ( clk, rst, A, B, product, overFlow );
  input [31:0] A;
  input [31:0] B;
  output [31:0] product;
  input clk, rst;
  output overFlow;
  wire   tempOverflow;
  wire   [31:0] in2;
  wire   [31:0] in1;
  wire   [31:0] out;

  DFF_X1 overFlow_reg ( .D(tempOverflow), .CK(clk), .Q(overFlow) );
  Register64bit inputRegister ( .clk(clk), .rst(rst), .in({B, A}), .out({in2, 
        in1}) );
  fpu fpua ( .in1(in1), .in2(in2), .overFlow(tempOverflow), .out(out) );
  Register32bit outRegister ( .clk(clk), .rst(rst), .in(out), .out(product) );
endmodule

